<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>12.8408,6.72322,152.792,-67.8785</PageViewport>
<gate>
<ID>2</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-17.5</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>55 </output>
<output>
<ID>OUT_1</ID>56 </output>
<output>
<ID>OUT_10</ID>65 </output>
<output>
<ID>OUT_11</ID>66 </output>
<output>
<ID>OUT_12</ID>67 </output>
<output>
<ID>OUT_13</ID>68 </output>
<output>
<ID>OUT_14</ID>69 </output>
<output>
<ID>OUT_15</ID>70 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>58 </output>
<output>
<ID>OUT_4</ID>59 </output>
<output>
<ID>OUT_5</ID>60 </output>
<output>
<ID>OUT_6</ID>61 </output>
<output>
<ID>OUT_7</ID>62 </output>
<output>
<ID>OUT_8</ID>63 </output>
<output>
<ID>OUT_9</ID>64 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>3</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-40.5</position>
<input>
<ID>ENABLE_0</ID>19 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>22 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_10</ID>44 </output>
<output>
<ID>OUT_11</ID>52 </output>
<output>
<ID>OUT_12</ID>45 </output>
<output>
<ID>OUT_13</ID>53 </output>
<output>
<ID>OUT_14</ID>46 </output>
<output>
<ID>OUT_15</ID>54 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>48 </output>
<output>
<ID>OUT_4</ID>41 </output>
<output>
<ID>OUT_5</ID>49 </output>
<output>
<ID>OUT_6</ID>42 </output>
<output>
<ID>OUT_7</ID>50 </output>
<output>
<ID>OUT_8</ID>43 </output>
<output>
<ID>OUT_9</ID>51 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>5</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>16 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-35</position>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>11 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>15 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-23</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>4 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>8 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-47</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>7 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>19.5,-36</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>19,-10</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>19,-22.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>19,-47.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BA_DECODER_2x4</type>
<position>60.5,-1</position>
<input>
<ID>ENABLE</ID>17 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>55.5,0.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>51,-2.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>56,3.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>44.5,-2</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-36.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>49 </input>
<input>
<ID>IN_3</ID>50 </input>
<input>
<ID>IN_B_0</ID>22 </input>
<input>
<ID>IN_B_1</ID>40 </input>
<input>
<ID>IN_B_2</ID>41 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<output>
<ID>carry_out</ID>21 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-52.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_B_0</ID>43 </input>
<input>
<ID>IN_B_1</ID>44 </input>
<input>
<ID>IN_B_2</ID>45 </input>
<input>
<ID>IN_B_3</ID>46 </input>
<output>
<ID>OUT_0</ID>75 </output>
<output>
<ID>OUT_1</ID>76 </output>
<output>
<ID>OUT_2</ID>77 </output>
<output>
<ID>OUT_3</ID>78 </output>
<input>
<ID>carry_in</ID>21 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>94,-29</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>94.5,-57.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>80,-30</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>80.5,-36.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>80,-46</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>81,-53</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>82,-26</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>87,-22.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>82,-19</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>87,-15.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>82,-12</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>87,-8.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>82,-5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>87,-1.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_MUX_2x1</type>
<position>112,-13</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>94 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_MUX_2x1</type>
<position>112,-18</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>93 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_MUX_2x1</type>
<position>112,-23</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>92 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_MUX_2x1</type>
<position>112,-28</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>91 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_MUX_2x1</type>
<position>112,-33</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>90 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_MUX_2x1</type>
<position>112,-38</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>112,-43</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>88 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_MUX_2x1</type>
<position>112,-48</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>87 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>134.5,-30</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>90 </input>
<input>
<ID>IN_4</ID>91 </input>
<input>
<ID>IN_5</ID>92 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>94 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 18</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>112,-51.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>113,-9</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>126,-40</position>
<input>
<ID>N_in2</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>128.5,-40</position>
<input>
<ID>N_in2</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>131,-40</position>
<input>
<ID>N_in2</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>133.5,-40</position>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>136,-40</position>
<input>
<ID>N_in2</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>138.5,-40</position>
<input>
<ID>N_in2</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>141,-40</position>
<input>
<ID>N_in2</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>143.5,-40</position>
<input>
<ID>N_in2</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>143.5,-42</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>141,-42</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>138.5,-42</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>136,-42</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>133.5,-42</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>131,-42</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>128.5,-42</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>126,-42</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-50,50.5,-48</points>
<intersection>-50 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-48,67,-48</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-50,50.5,-50</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-48,67,-25</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-47,50.5,-24</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection>
<intersection>-24 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-47,67,-47</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-26,50.5,-26</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-24,67,-24</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-48,50.5,-46</points>
<intersection>-48 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-46,67,-46</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-48,50.5,-48</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-46,67,-23</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-45,50.5,-22</points>
<intersection>-45 1</intersection>
<intersection>-24 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-45,67,-45</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-24,50.5,-24</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-22,67,-22</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-46,50.5,-44</points>
<intersection>-46 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-44,67,-44</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-46,50.5,-46</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-44,67,-21</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-43,50.5,-20</points>
<intersection>-43 1</intersection>
<intersection>-22 2</intersection>
<intersection>-20 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-43,67,-43</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-22,50.5,-22</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-20,67,-20</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-44,50.5,-42</points>
<intersection>-44 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-42,67,-42</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-44,50.5,-44</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-42,67,-19</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-41,50.5,-18</points>
<intersection>-41 1</intersection>
<intersection>-20 2</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-41,67,-41</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-20,50.5,-20</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-18,67,-18</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-40,50.5,-17</points>
<intersection>-40 1</intersection>
<intersection>-38 2</intersection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-40,67,-40</points>
<connection>
<GID>3</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-38,50.5,-38</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-17,67,-17</points>
<connection>
<GID>2</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-39,50.5,-14</points>
<intersection>-39 1</intersection>
<intersection>-16 4</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-39,67,-39</points>
<connection>
<GID>3</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-14,50.5,-14</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-16,67,-16</points>
<connection>
<GID>2</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-38,50.5,-15</points>
<intersection>-38 1</intersection>
<intersection>-36 2</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-38,67,-38</points>
<connection>
<GID>3</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-36,50.5,-36</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-15,67,-15</points>
<connection>
<GID>2</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-37,50.5,-12</points>
<intersection>-37 1</intersection>
<intersection>-14 3</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-37,67,-37</points>
<connection>
<GID>3</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-12,50.5,-12</points>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-14,67,-14</points>
<connection>
<GID>2</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-36,50.5,-13</points>
<intersection>-36 1</intersection>
<intersection>-34 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-36,67,-36</points>
<connection>
<GID>3</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-34,50.5,-34</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-13,67,-13</points>
<connection>
<GID>2</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-35,50.5,-10</points>
<intersection>-35 1</intersection>
<intersection>-12 3</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-35,67,-35</points>
<connection>
<GID>3</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-10,50.5,-10</points>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-12,67,-12</points>
<connection>
<GID>2</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-34,50.5,-11</points>
<intersection>-34 1</intersection>
<intersection>-32 2</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-34,67,-34</points>
<connection>
<GID>3</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-32,50.5,-32</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-11,67,-11</points>
<connection>
<GID>2</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-33,50.5,-8</points>
<intersection>-33 1</intersection>
<intersection>-10 3</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-33,67,-33</points>
<connection>
<GID>3</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-8,50.5,-8</points>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-10,67,-10</points>
<connection>
<GID>2</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,0.5,57.5,0.5</points>
<connection>
<GID>15</GID>
<name>ENABLE</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,6,109,6</points>
<intersection>53 8</intersection>
<intersection>109 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>109,-45.5,109,6</points>
<intersection>-45.5 18</intersection>
<intersection>-40.5 19</intersection>
<intersection>-35.5 20</intersection>
<intersection>-30.5 21</intersection>
<intersection>-25.5 22</intersection>
<intersection>-20.5 23</intersection>
<intersection>-15.5 24</intersection>
<intersection>-10.5 25</intersection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>53,-2.5,53,6</points>
<intersection>-2.5 10</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>53,-2.5,57.5,-2.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>53 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>109,-45.5,112,-45.5</points>
<connection>
<GID>54</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>109,-40.5,112,-40.5</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>109,-35.5,112,-35.5</points>
<connection>
<GID>52</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>109,-30.5,112,-30.5</points>
<connection>
<GID>51</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>109,-25.5,112,-25.5</points>
<connection>
<GID>50</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>109,-20.5,112,-20.5</points>
<connection>
<GID>49</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>109,-15.5,112,-15.5</points>
<connection>
<GID>48</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>109,-10.5,112,-10.5</points>
<connection>
<GID>47</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-31.5,64.5,-2.5</points>
<intersection>-31.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-2.5,64.5,-2.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-31.5,69,-31.5</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-8.5,69,-1.5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-1.5,69,-1.5</points>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-44.5,85.5,-44.5</points>
<connection>
<GID>25</GID>
<name>carry_out</name></connection>
<connection>
<GID>26</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-48,72.5,-31.5</points>
<intersection>-48 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-31.5,82.5,-31.5</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-48,72.5,-48</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-46,73,-32.5</points>
<intersection>-46 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-32.5,82.5,-32.5</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-46,73,-46</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-44,73.5,-33.5</points>
<intersection>-44 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-33.5,82.5,-33.5</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-44,73.5,-44</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-42,74,-34.5</points>
<intersection>-42 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-34.5,82.5,-34.5</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-42,74,-42</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-47.5,76,-40</points>
<intersection>-47.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-47.5,82.5,-47.5</points>
<connection>
<GID>26</GID>
<name>IN_B_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-40,76,-40</points>
<connection>
<GID>3</GID>
<name>OUT_8</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-48.5,75.5,-38</points>
<intersection>-48.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-48.5,82.5,-48.5</points>
<connection>
<GID>26</GID>
<name>IN_B_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-38,75.5,-38</points>
<connection>
<GID>3</GID>
<name>OUT_10</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-49.5,75,-36</points>
<intersection>-49.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-49.5,82.5,-49.5</points>
<connection>
<GID>26</GID>
<name>IN_B_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-36,75,-36</points>
<connection>
<GID>3</GID>
<name>OUT_12</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-50.5,74.5,-34</points>
<intersection>-50.5 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-50.5,82.5,-50.5</points>
<connection>
<GID>26</GID>
<name>IN_B_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-34,74.5,-34</points>
<connection>
<GID>3</GID>
<name>OUT_14</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-47,76.5,-38.5</points>
<intersection>-47 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-38.5,82.5,-38.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-47,76.5,-47</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-45,76.5,-39.5</points>
<intersection>-45 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-39.5,82.5,-39.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-45,76.5,-45</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-43,76.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-40.5,82.5,-40.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-43,76.5,-43</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-41.5,76.5,-41</points>
<intersection>-41.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-41.5,82.5,-41.5</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-41,76.5,-41</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-54.5,78.5,-39</points>
<intersection>-54.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-54.5,82.5,-54.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-39,78.5,-39</points>
<connection>
<GID>3</GID>
<name>OUT_9</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-55.5,78,-37</points>
<intersection>-55.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-55.5,82.5,-55.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-37,78,-37</points>
<connection>
<GID>3</GID>
<name>OUT_11</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-56.5,77.5,-35</points>
<intersection>-56.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-56.5,82.5,-56.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-35,77.5,-35</points>
<connection>
<GID>3</GID>
<name>OUT_13</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-57.5,77,-33</points>
<intersection>-57.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-57.5,82.5,-57.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-33,77,-33</points>
<connection>
<GID>3</GID>
<name>OUT_15</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-27,72,-25</points>
<intersection>-27 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-27,79,-27</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-25,72,-25</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-25,79,-25</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-25,71,-24</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-23.5,74.5,-23</points>
<intersection>-23.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-23.5,84,-23.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-23,74.5,-23</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-21.5,84,-21.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-22,71,-21.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-20,79,-20</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-21,71,-20</points>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-20,72,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-18,79,-18</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-20,72,-20</points>
<connection>
<GID>2</GID>
<name>OUT_5</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-19,73,-16.5</points>
<intersection>-19 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-16.5,84,-16.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-19,73,-19</points>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-18,72.5,-14.5</points>
<intersection>-18 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-14.5,84,-14.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-18,72.5,-18</points>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-17,72,-13</points>
<intersection>-17 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-13,79,-13</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-17,72,-17</points>
<connection>
<GID>2</GID>
<name>OUT_8</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-16,72,-11</points>
<intersection>-16 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-11,79,-11</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-16,72,-16</points>
<connection>
<GID>2</GID>
<name>OUT_9</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-15,72.5,-9.5</points>
<intersection>-15 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-9.5,84,-9.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-15,72.5,-15</points>
<connection>
<GID>2</GID>
<name>OUT_10</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-14,72.5,-7.5</points>
<intersection>-14 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-7.5,84,-7.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-14,72.5,-14</points>
<connection>
<GID>2</GID>
<name>OUT_11</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-13,72,-6</points>
<intersection>-13 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-6,79,-6</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-13,72,-13</points>
<connection>
<GID>2</GID>
<name>OUT_12</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-12,72,-4</points>
<intersection>-12 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4,79,-4</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-12,72,-12</points>
<connection>
<GID>2</GID>
<name>OUT_13</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-11,71.5,-2.5</points>
<intersection>-11 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-2.5,84,-2.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-11,71.5,-11</points>
<connection>
<GID>2</GID>
<name>OUT_14</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-10,71,-0.5</points>
<connection>
<GID>2</GID>
<name>OUT_15</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-0.5,84,-0.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-49,100,-35</points>
<intersection>-49 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-49,110,-49</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-35,100,-35</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-44,100,-36</points>
<intersection>-44 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-44,110,-44</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-36,100,-36</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-39,100,-37</points>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-39,110,-39</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-37,100,-37</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-38,100,-34</points>
<intersection>-38 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-34,110,-34</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-38,100,-38</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-51,100,-29</points>
<intersection>-51 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-29,110,-29</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-51,100,-51</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-52,100,-24</points>
<intersection>-52 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-24,110,-24</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-52,100,-52</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-53,100,-19</points>
<intersection>-53 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-19,110,-19</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-53,100,-53</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-54,100,-14</points>
<intersection>-54 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-14,110,-14</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-54,100,-54</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-47,97.5,-26</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-47,110,-47</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-26,97.5,-26</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-42,100,-22.5</points>
<intersection>-42 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-22.5,100,-22.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-42,110,-42</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-37,97.5,-19</points>
<intersection>-37 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-19,97.5,-19</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-37,110,-37</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-32,100,-15.5</points>
<intersection>-32 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-15.5,100,-15.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-32,110,-32</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-27,97.5,-12</points>
<intersection>-27 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-12,97.5,-12</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-27,110,-27</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-22,100,-8.5</points>
<intersection>-22 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-8.5,100,-8.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-22,110,-22</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-17,97.5,-5</points>
<intersection>-17 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-5,97.5,-5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-17,110,-17</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-12,100,-1.5</points>
<intersection>-12 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-1.5,100,-1.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-12,110,-12</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-48,121.5,-33</points>
<intersection>-48 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-33,129.5,-33</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection>
<intersection>122.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-48,121.5,-48</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>122.5,-38.5,122.5,-33</points>
<intersection>-38.5 8</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-38.5,143.5,-38.5</points>
<intersection>122.5 7</intersection>
<intersection>143.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>143.5,-39,143.5,-38.5</points>
<connection>
<GID>86</GID>
<name>N_in2</name></connection>
<intersection>-38.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-43,121.5,-32</points>
<intersection>-43 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-32,129.5,-32</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection>
<intersection>123 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-43,121.5,-43</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123,-38,123,-32</points>
<intersection>-38 8</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123,-38,141,-38</points>
<intersection>123 7</intersection>
<intersection>141 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>141,-39,141,-38</points>
<connection>
<GID>85</GID>
<name>N_in2</name></connection>
<intersection>-38 8</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-38,121.5,-31</points>
<intersection>-38 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-31,129.5,-31</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>121.5 0</intersection>
<intersection>123.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-38,121.5,-38</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123.5,-37.5,123.5,-31</points>
<intersection>-37.5 8</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123.5,-37.5,138.5,-37.5</points>
<intersection>123.5 7</intersection>
<intersection>138.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>138.5,-39,138.5,-37.5</points>
<connection>
<GID>84</GID>
<name>N_in2</name></connection>
<intersection>-37.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-33,121.5,-30</points>
<intersection>-33 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-30,129.5,-30</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>121.5 0</intersection>
<intersection>124 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-33,121.5,-33</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124,-37,124,-30</points>
<intersection>-37 9</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124,-37,136,-37</points>
<intersection>124 8</intersection>
<intersection>136 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>136,-39,136,-37</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>-37 9</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-29,121.5,-28</points>
<intersection>-29 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-29,129.5,-29</points>
<connection>
<GID>56</GID>
<name>IN_4</name></connection>
<intersection>121.5 0</intersection>
<intersection>124.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-28,121.5,-28</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124.5,-36.5,124.5,-29</points>
<intersection>-36.5 9</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124.5,-36.5,133.5,-36.5</points>
<intersection>124.5 8</intersection>
<intersection>133.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>133.5,-39,133.5,-36.5</points>
<connection>
<GID>82</GID>
<name>N_in2</name></connection>
<intersection>-36.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-28,121.5,-23</points>
<intersection>-28 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-28,129.5,-28</points>
<connection>
<GID>56</GID>
<name>IN_5</name></connection>
<intersection>121.5 0</intersection>
<intersection>125 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-23,121.5,-23</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125,-36,125,-28</points>
<intersection>-36 8</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125,-36,131,-36</points>
<intersection>125 7</intersection>
<intersection>131 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>131,-39,131,-36</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<intersection>-36 8</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-27,121.5,-18</points>
<intersection>-27 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-27,129.5,-27</points>
<connection>
<GID>56</GID>
<name>IN_6</name></connection>
<intersection>121.5 0</intersection>
<intersection>125.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-18,121.5,-18</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125.5,-35.5,125.5,-27</points>
<intersection>-35.5 8</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125.5,-35.5,128.5,-35.5</points>
<intersection>125.5 7</intersection>
<intersection>128.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>128.5,-39,128.5,-35.5</points>
<connection>
<GID>80</GID>
<name>N_in2</name></connection>
<intersection>-35.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-26,121.5,-13</points>
<intersection>-26 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-13,121.5,-13</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-26,129.5,-26</points>
<connection>
<GID>56</GID>
<name>IN_7</name></connection>
<intersection>121.5 0</intersection>
<intersection>126 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>126,-39,126,-26</points>
<connection>
<GID>79</GID>
<name>N_in2</name></connection>
<intersection>-26 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 1>
<page 2>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 2>
<page 3>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 3>
<page 4>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 4>
<page 5>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 5>
<page 6>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 6>
<page 7>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 7>
<page 8>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 8>
<page 9>
<PageViewport>0,0.364097,146.309,-77.6262</PageViewport></page 9></circuit>