<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.25,40.8679,539.303,-229.927</PageViewport>
<gate>
<ID>2</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-17.5</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>55 </output>
<output>
<ID>OUT_1</ID>56 </output>
<output>
<ID>OUT_10</ID>65 </output>
<output>
<ID>OUT_11</ID>66 </output>
<output>
<ID>OUT_12</ID>67 </output>
<output>
<ID>OUT_13</ID>68 </output>
<output>
<ID>OUT_14</ID>69 </output>
<output>
<ID>OUT_15</ID>70 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>58 </output>
<output>
<ID>OUT_4</ID>59 </output>
<output>
<ID>OUT_5</ID>60 </output>
<output>
<ID>OUT_6</ID>61 </output>
<output>
<ID>OUT_7</ID>62 </output>
<output>
<ID>OUT_8</ID>63 </output>
<output>
<ID>OUT_9</ID>64 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>3</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-40.5</position>
<input>
<ID>ENABLE_0</ID>19 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>22 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_10</ID>44 </output>
<output>
<ID>OUT_11</ID>52 </output>
<output>
<ID>OUT_12</ID>45 </output>
<output>
<ID>OUT_13</ID>53 </output>
<output>
<ID>OUT_14</ID>46 </output>
<output>
<ID>OUT_15</ID>54 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>48 </output>
<output>
<ID>OUT_4</ID>41 </output>
<output>
<ID>OUT_5</ID>49 </output>
<output>
<ID>OUT_6</ID>42 </output>
<output>
<ID>OUT_7</ID>50 </output>
<output>
<ID>OUT_8</ID>43 </output>
<output>
<ID>OUT_9</ID>51 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>46.5,-4.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>16 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-35</position>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>11 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>15 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>7</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-23</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>4 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>8 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-47</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>7 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>19.5,-36</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>19,-10</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>19,-22.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>19,-47.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BA_DECODER_2x4</type>
<position>60.5,-1</position>
<input>
<ID>ENABLE</ID>17 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>55.5,0.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>51,-2.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>56,3.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>44.5,-2</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-36.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>49 </input>
<input>
<ID>IN_3</ID>50 </input>
<input>
<ID>IN_B_0</ID>22 </input>
<input>
<ID>IN_B_1</ID>40 </input>
<input>
<ID>IN_B_2</ID>41 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<output>
<ID>carry_out</ID>21 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-52.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_B_0</ID>43 </input>
<input>
<ID>IN_B_1</ID>44 </input>
<input>
<ID>IN_B_2</ID>45 </input>
<input>
<ID>IN_B_3</ID>46 </input>
<output>
<ID>OUT_0</ID>75 </output>
<output>
<ID>OUT_1</ID>76 </output>
<output>
<ID>OUT_2</ID>77 </output>
<output>
<ID>OUT_3</ID>78 </output>
<input>
<ID>carry_in</ID>21 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>94,-29</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>94.5,-57.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>80,-30</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>80.5,-36.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>80,-46</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>81,-53</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>82,-26</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>87,-22.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>82,-19</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>87,-15.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>82,-12</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>87,-8.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>82,-5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>87,-1.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_MUX_2x1</type>
<position>112,-13</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>94 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_MUX_2x1</type>
<position>112,-18</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>93 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_MUX_2x1</type>
<position>112,-23</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>92 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_MUX_2x1</type>
<position>112,-28</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>91 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_MUX_2x1</type>
<position>112,-33</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>90 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_MUX_2x1</type>
<position>112,-38</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>112,-43</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>88 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_MUX_2x1</type>
<position>112,-48</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>87 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>134.5,-30</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>90 </input>
<input>
<ID>IN_4</ID>91 </input>
<input>
<ID>IN_5</ID>92 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>94 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>112,-51.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>113,-9</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>126,-40</position>
<input>
<ID>N_in2</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>128.5,-40</position>
<input>
<ID>N_in2</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>131,-40</position>
<input>
<ID>N_in2</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>133.5,-40</position>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>136,-40</position>
<input>
<ID>N_in2</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>138.5,-40</position>
<input>
<ID>N_in2</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>141,-40</position>
<input>
<ID>N_in2</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>143.5,-40</position>
<input>
<ID>N_in2</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>143.5,-42</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>141,-42</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>138.5,-42</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>136,-42</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>133.5,-42</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>131,-42</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>128.5,-42</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>126,-42</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-50,50.5,-48</points>
<intersection>-50 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-48,67,-48</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-50,50.5,-50</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-48,67,-25</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-47,50.5,-24</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection>
<intersection>-24 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-47,67,-47</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-26,50.5,-26</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-24,67,-24</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-48,50.5,-46</points>
<intersection>-48 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-46,67,-46</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-48,50.5,-48</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-46,67,-23</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-45,50.5,-22</points>
<intersection>-45 1</intersection>
<intersection>-24 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-45,67,-45</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-24,50.5,-24</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-22,67,-22</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-46,50.5,-44</points>
<intersection>-46 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-44,67,-44</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-46,50.5,-46</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-44,67,-21</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-43,50.5,-20</points>
<intersection>-43 1</intersection>
<intersection>-22 2</intersection>
<intersection>-20 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-43,67,-43</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-22,50.5,-22</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-20,67,-20</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-44,50.5,-42</points>
<intersection>-44 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-42,67,-42</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-44,50.5,-44</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-42,67,-19</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-41,50.5,-18</points>
<intersection>-41 1</intersection>
<intersection>-20 2</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-41,67,-41</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-20,50.5,-20</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-18,67,-18</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-40,50.5,-17</points>
<intersection>-40 1</intersection>
<intersection>-38 2</intersection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-40,67,-40</points>
<connection>
<GID>3</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-38,50.5,-38</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-17,67,-17</points>
<connection>
<GID>2</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-39,50.5,-14</points>
<intersection>-39 1</intersection>
<intersection>-16 4</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-39,67,-39</points>
<connection>
<GID>3</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-14,50.5,-14</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-16,67,-16</points>
<connection>
<GID>2</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-38,50.5,-15</points>
<intersection>-38 1</intersection>
<intersection>-36 2</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-38,67,-38</points>
<connection>
<GID>3</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-36,50.5,-36</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-15,67,-15</points>
<connection>
<GID>2</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-37,50.5,-12</points>
<intersection>-37 1</intersection>
<intersection>-14 3</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-37,67,-37</points>
<connection>
<GID>3</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-12,50.5,-12</points>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-14,67,-14</points>
<connection>
<GID>2</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-36,50.5,-13</points>
<intersection>-36 1</intersection>
<intersection>-34 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-36,67,-36</points>
<connection>
<GID>3</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-34,50.5,-34</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-13,67,-13</points>
<connection>
<GID>2</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-35,50.5,-10</points>
<intersection>-35 1</intersection>
<intersection>-12 3</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-35,67,-35</points>
<connection>
<GID>3</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-10,50.5,-10</points>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-12,67,-12</points>
<connection>
<GID>2</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-34,50.5,-11</points>
<intersection>-34 1</intersection>
<intersection>-32 2</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-34,67,-34</points>
<connection>
<GID>3</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-32,50.5,-32</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-11,67,-11</points>
<connection>
<GID>2</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-33,50.5,-8</points>
<intersection>-33 1</intersection>
<intersection>-10 3</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-33,67,-33</points>
<connection>
<GID>3</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-8,50.5,-8</points>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-10,67,-10</points>
<connection>
<GID>2</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,0.5,57.5,0.5</points>
<connection>
<GID>15</GID>
<name>ENABLE</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,6,109,6</points>
<intersection>53 8</intersection>
<intersection>109 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>109,-45.5,109,6</points>
<intersection>-45.5 18</intersection>
<intersection>-40.5 19</intersection>
<intersection>-35.5 20</intersection>
<intersection>-30.5 21</intersection>
<intersection>-25.5 22</intersection>
<intersection>-20.5 23</intersection>
<intersection>-15.5 24</intersection>
<intersection>-10.5 25</intersection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>53,-2.5,53,6</points>
<intersection>-2.5 10</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>53,-2.5,57.5,-2.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>53 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>109,-45.5,112,-45.5</points>
<connection>
<GID>54</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>109,-40.5,112,-40.5</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>109,-35.5,112,-35.5</points>
<connection>
<GID>52</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>109,-30.5,112,-30.5</points>
<connection>
<GID>51</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>109,-25.5,112,-25.5</points>
<connection>
<GID>50</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>109,-20.5,112,-20.5</points>
<connection>
<GID>49</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>109,-15.5,112,-15.5</points>
<connection>
<GID>48</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>109,-10.5,112,-10.5</points>
<connection>
<GID>47</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-31.5,64.5,-2.5</points>
<intersection>-31.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-2.5,64.5,-2.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-31.5,69,-31.5</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-8.5,69,-1.5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-1.5,69,-1.5</points>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-44.5,85.5,-44.5</points>
<connection>
<GID>25</GID>
<name>carry_out</name></connection>
<connection>
<GID>26</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-48,72.5,-31.5</points>
<intersection>-48 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-31.5,82.5,-31.5</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-48,72.5,-48</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-46,73,-32.5</points>
<intersection>-46 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-32.5,82.5,-32.5</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-46,73,-46</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-44,73.5,-33.5</points>
<intersection>-44 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-33.5,82.5,-33.5</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-44,73.5,-44</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-42,74,-34.5</points>
<intersection>-42 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-34.5,82.5,-34.5</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-42,74,-42</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-47.5,76,-40</points>
<intersection>-47.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-47.5,82.5,-47.5</points>
<connection>
<GID>26</GID>
<name>IN_B_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-40,76,-40</points>
<connection>
<GID>3</GID>
<name>OUT_8</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-48.5,75.5,-38</points>
<intersection>-48.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-48.5,82.5,-48.5</points>
<connection>
<GID>26</GID>
<name>IN_B_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-38,75.5,-38</points>
<connection>
<GID>3</GID>
<name>OUT_10</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-49.5,75,-36</points>
<intersection>-49.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-49.5,82.5,-49.5</points>
<connection>
<GID>26</GID>
<name>IN_B_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-36,75,-36</points>
<connection>
<GID>3</GID>
<name>OUT_12</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-50.5,74.5,-34</points>
<intersection>-50.5 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-50.5,82.5,-50.5</points>
<connection>
<GID>26</GID>
<name>IN_B_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-34,74.5,-34</points>
<connection>
<GID>3</GID>
<name>OUT_14</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-47,76.5,-38.5</points>
<intersection>-47 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-38.5,82.5,-38.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-47,76.5,-47</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-45,76.5,-39.5</points>
<intersection>-45 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-39.5,82.5,-39.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-45,76.5,-45</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-43,76.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-40.5,82.5,-40.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-43,76.5,-43</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-41.5,76.5,-41</points>
<intersection>-41.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-41.5,82.5,-41.5</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-41,76.5,-41</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-54.5,78.5,-39</points>
<intersection>-54.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-54.5,82.5,-54.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-39,78.5,-39</points>
<connection>
<GID>3</GID>
<name>OUT_9</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-55.5,78,-37</points>
<intersection>-55.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-55.5,82.5,-55.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-37,78,-37</points>
<connection>
<GID>3</GID>
<name>OUT_11</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-56.5,77.5,-35</points>
<intersection>-56.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-56.5,82.5,-56.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-35,77.5,-35</points>
<connection>
<GID>3</GID>
<name>OUT_13</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-57.5,77,-33</points>
<intersection>-57.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-57.5,82.5,-57.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-33,77,-33</points>
<connection>
<GID>3</GID>
<name>OUT_15</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-27,72,-25</points>
<intersection>-27 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-27,79,-27</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-25,72,-25</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-25,79,-25</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-25,71,-24</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-23.5,74.5,-23</points>
<intersection>-23.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-23.5,84,-23.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-23,74.5,-23</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-21.5,84,-21.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-22,71,-21.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-20,79,-20</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-21,71,-20</points>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-20,72,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-18,79,-18</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-20,72,-20</points>
<connection>
<GID>2</GID>
<name>OUT_5</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-19,73,-16.5</points>
<intersection>-19 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-16.5,84,-16.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-19,73,-19</points>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-18,72.5,-14.5</points>
<intersection>-18 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-14.5,84,-14.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-18,72.5,-18</points>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-17,72,-13</points>
<intersection>-17 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-13,79,-13</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-17,72,-17</points>
<connection>
<GID>2</GID>
<name>OUT_8</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-16,72,-11</points>
<intersection>-16 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-11,79,-11</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-16,72,-16</points>
<connection>
<GID>2</GID>
<name>OUT_9</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-15,72.5,-9.5</points>
<intersection>-15 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-9.5,84,-9.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-15,72.5,-15</points>
<connection>
<GID>2</GID>
<name>OUT_10</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-14,72.5,-7.5</points>
<intersection>-14 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-7.5,84,-7.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-14,72.5,-14</points>
<connection>
<GID>2</GID>
<name>OUT_11</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-13,72,-6</points>
<intersection>-13 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-6,79,-6</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-13,72,-13</points>
<connection>
<GID>2</GID>
<name>OUT_12</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-12,72,-4</points>
<intersection>-12 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4,79,-4</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-12,72,-12</points>
<connection>
<GID>2</GID>
<name>OUT_13</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-11,71.5,-2.5</points>
<intersection>-11 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-2.5,84,-2.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-11,71.5,-11</points>
<connection>
<GID>2</GID>
<name>OUT_14</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-10,71,-0.5</points>
<connection>
<GID>2</GID>
<name>OUT_15</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-0.5,84,-0.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-49,100,-35</points>
<intersection>-49 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-49,110,-49</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-35,100,-35</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-44,100,-36</points>
<intersection>-44 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-44,110,-44</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-36,100,-36</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-39,100,-37</points>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-39,110,-39</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-37,100,-37</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-38,100,-34</points>
<intersection>-38 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-34,110,-34</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-38,100,-38</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-51,100,-29</points>
<intersection>-51 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-29,110,-29</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-51,100,-51</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-52,100,-24</points>
<intersection>-52 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-24,110,-24</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-52,100,-52</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-53,100,-19</points>
<intersection>-53 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-19,110,-19</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-53,100,-53</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-54,100,-14</points>
<intersection>-54 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-14,110,-14</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-54,100,-54</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-47,97.5,-26</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-47,110,-47</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-26,97.5,-26</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-42,100,-22.5</points>
<intersection>-42 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-22.5,100,-22.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-42,110,-42</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-37,97.5,-19</points>
<intersection>-37 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-19,97.5,-19</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-37,110,-37</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-32,100,-15.5</points>
<intersection>-32 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-15.5,100,-15.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-32,110,-32</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-27,97.5,-12</points>
<intersection>-27 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-12,97.5,-12</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-27,110,-27</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-22,100,-8.5</points>
<intersection>-22 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-8.5,100,-8.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-22,110,-22</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-17,97.5,-5</points>
<intersection>-17 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-5,97.5,-5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-17,110,-17</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-12,100,-1.5</points>
<intersection>-12 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-1.5,100,-1.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-12,110,-12</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-48,121.5,-33</points>
<intersection>-48 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-33,129.5,-33</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection>
<intersection>122.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-48,121.5,-48</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>122.5,-38.5,122.5,-33</points>
<intersection>-38.5 8</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-38.5,143.5,-38.5</points>
<intersection>122.5 7</intersection>
<intersection>143.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>143.5,-39,143.5,-38.5</points>
<connection>
<GID>86</GID>
<name>N_in2</name></connection>
<intersection>-38.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-43,121.5,-32</points>
<intersection>-43 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-32,129.5,-32</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection>
<intersection>123 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-43,121.5,-43</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123,-38,123,-32</points>
<intersection>-38 8</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123,-38,141,-38</points>
<intersection>123 7</intersection>
<intersection>141 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>141,-39,141,-38</points>
<connection>
<GID>85</GID>
<name>N_in2</name></connection>
<intersection>-38 8</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-38,121.5,-31</points>
<intersection>-38 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-31,129.5,-31</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>121.5 0</intersection>
<intersection>123.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-38,121.5,-38</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123.5,-37.5,123.5,-31</points>
<intersection>-37.5 8</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123.5,-37.5,138.5,-37.5</points>
<intersection>123.5 7</intersection>
<intersection>138.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>138.5,-39,138.5,-37.5</points>
<connection>
<GID>84</GID>
<name>N_in2</name></connection>
<intersection>-37.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-33,121.5,-30</points>
<intersection>-33 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-30,129.5,-30</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>121.5 0</intersection>
<intersection>124 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-33,121.5,-33</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124,-37,124,-30</points>
<intersection>-37 9</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124,-37,136,-37</points>
<intersection>124 8</intersection>
<intersection>136 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>136,-39,136,-37</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>-37 9</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-29,121.5,-28</points>
<intersection>-29 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-29,129.5,-29</points>
<connection>
<GID>56</GID>
<name>IN_4</name></connection>
<intersection>121.5 0</intersection>
<intersection>124.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-28,121.5,-28</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124.5,-36.5,124.5,-29</points>
<intersection>-36.5 9</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124.5,-36.5,133.5,-36.5</points>
<intersection>124.5 8</intersection>
<intersection>133.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>133.5,-39,133.5,-36.5</points>
<connection>
<GID>82</GID>
<name>N_in2</name></connection>
<intersection>-36.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-28,121.5,-23</points>
<intersection>-28 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-28,129.5,-28</points>
<connection>
<GID>56</GID>
<name>IN_5</name></connection>
<intersection>121.5 0</intersection>
<intersection>125 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-23,121.5,-23</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125,-36,125,-28</points>
<intersection>-36 8</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125,-36,131,-36</points>
<intersection>125 7</intersection>
<intersection>131 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>131,-39,131,-36</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<intersection>-36 8</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-27,121.5,-18</points>
<intersection>-27 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-27,129.5,-27</points>
<connection>
<GID>56</GID>
<name>IN_6</name></connection>
<intersection>121.5 0</intersection>
<intersection>125.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-18,121.5,-18</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125.5,-35.5,125.5,-27</points>
<intersection>-35.5 8</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125.5,-35.5,128.5,-35.5</points>
<intersection>125.5 7</intersection>
<intersection>128.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>128.5,-39,128.5,-35.5</points>
<connection>
<GID>80</GID>
<name>N_in2</name></connection>
<intersection>-35.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-26,121.5,-13</points>
<intersection>-26 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-13,121.5,-13</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-26,129.5,-26</points>
<connection>
<GID>56</GID>
<name>IN_7</name></connection>
<intersection>121.5 0</intersection>
<intersection>126 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>126,-39,126,-26</points>
<connection>
<GID>79</GID>
<name>N_in2</name></connection>
<intersection>-26 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-27.5273,337.155,1750.47,-579.844</PageViewport>
<gate>
<ID>1</ID>
<type>AE_RAM_8x8</type>
<position>59.5,-99.5</position>
<input>
<ID>ADDRESS_0</ID>98 </input>
<input>
<ID>ADDRESS_1</ID>102 </input>
<input>
<ID>ADDRESS_2</ID>97 </input>
<input>
<ID>ADDRESS_3</ID>100 </input>
<input>
<ID>ADDRESS_4</ID>99 </input>
<input>
<ID>ADDRESS_5</ID>101 </input>
<input>
<ID>ADDRESS_6</ID>103 </input>
<input>
<ID>ADDRESS_7</ID>96 </input>
<input>
<ID>DATA_IN_0</ID>25 </input>
<input>
<ID>DATA_IN_1</ID>26 </input>
<input>
<ID>DATA_IN_2</ID>27 </input>
<input>
<ID>DATA_IN_3</ID>28 </input>
<input>
<ID>DATA_IN_4</ID>29 </input>
<input>
<ID>DATA_IN_5</ID>30 </input>
<input>
<ID>DATA_IN_6</ID>31 </input>
<input>
<ID>DATA_IN_7</ID>32 </input>
<output>
<ID>DATA_OUT_0</ID>25 </output>
<output>
<ID>DATA_OUT_1</ID>26 </output>
<output>
<ID>DATA_OUT_2</ID>27 </output>
<output>
<ID>DATA_OUT_3</ID>28 </output>
<output>
<ID>DATA_OUT_4</ID>29 </output>
<output>
<ID>DATA_OUT_5</ID>30 </output>
<output>
<ID>DATA_OUT_6</ID>31 </output>
<output>
<ID>DATA_OUT_7</ID>32 </output>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>write_clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>9</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>66,-113</position>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>28 </input>
<input>
<ID>IN_4</ID>29 </input>
<input>
<ID>IN_5</ID>30 </input>
<input>
<ID>IN_6</ID>31 </input>
<input>
<ID>IN_7</ID>32 </input>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>34 </output>
<output>
<ID>OUT_2</ID>35 </output>
<output>
<ID>OUT_3</ID>36 </output>
<output>
<ID>OUT_4</ID>37 </output>
<output>
<ID>OUT_5</ID>38 </output>
<output>
<ID>OUT_6</ID>39 </output>
<output>
<ID>OUT_7</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>14</ID>
<type>EE_VDD</type>
<position>67,-100</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>BB_CLOCK</type>
<position>24,-91.5</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>70.5,-113</position>
<input>
<ID>N_in0</ID>95 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>72.5,-113</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>74.5,-113</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>76.5,-113</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>78.5,-113</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>166.5,-34</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>80.5,-113</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>82.5,-113</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>166.5,-45</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>84.5,-113</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AE_REGISTER8</type>
<position>41,-100</position>
<output>
<ID>OUT_0</ID>98 </output>
<output>
<ID>OUT_1</ID>102 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>100 </output>
<output>
<ID>OUT_4</ID>99 </output>
<output>
<ID>OUT_5</ID>101 </output>
<output>
<ID>OUT_6</ID>103 </output>
<output>
<ID>OUT_7</ID>96 </output>
<input>
<ID>clock</ID>104 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_MUX_2x1</type>
<position>30,-108</position>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AE_REGISTER8</type>
<position>109.5,-45</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>128 </output>
<output>
<ID>OUT_1</ID>127 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>125 </output>
<output>
<ID>OUT_4</ID>124 </output>
<output>
<ID>OUT_5</ID>123 </output>
<output>
<ID>OUT_6</ID>122 </output>
<output>
<ID>OUT_7</ID>121 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>168 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_REGISTER8</type>
<position>109.5,-58</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>144 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>133 </output>
<output>
<ID>OUT_4</ID>132 </output>
<output>
<ID>OUT_5</ID>131 </output>
<output>
<ID>OUT_6</ID>130 </output>
<output>
<ID>OUT_7</ID>129 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>169 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_MUX_4x1</type>
<position>135,-7.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>136 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_MUX_4x1</type>
<position>135,-18.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>122 </input>
<input>
<ID>IN_2</ID>114 </input>
<input>
<ID>IN_3</ID>106 </input>
<output>
<ID>OUT</ID>137 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_MUX_4x1</type>
<position>135,-29.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT</ID>138 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_MUX_4x1</type>
<position>135,-39</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>108 </input>
<output>
<ID>OUT</ID>139 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_MUX_4x1</type>
<position>135,-50</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>117 </input>
<input>
<ID>IN_3</ID>109 </input>
<output>
<ID>OUT</ID>140 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_MUX_4x1</type>
<position>135,-61</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_MUX_4x1</type>
<position>135,-71.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>119 </input>
<input>
<ID>IN_3</ID>111 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_MUX_4x1</type>
<position>135,-82.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>112 </input>
<output>
<ID>OUT</ID>143 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>167,-40</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>140 </input>
<input>
<ID>IN_4</ID>139 </input>
<input>
<ID>IN_5</ID>138 </input>
<input>
<ID>IN_6</ID>137 </input>
<input>
<ID>IN_7</ID>136 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>71</ID>
<type>DD_KEYPAD_HEX</type>
<position>76.5,-22.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<output>
<ID>OUT_1</ID>147 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>BB_CLOCK</type>
<position>98,-66.5</position>
<output>
<ID>CLK</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>110.5,-11.5</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>110.5,-24.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>110.5,-38</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>110.5,-51</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>75,-15.5</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>DD_KEYPAD_HEX</type>
<position>76.5,-36.5</position>
<output>
<ID>OUT_0</ID>156 </output>
<output>
<ID>OUT_1</ID>157 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-7.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>148 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-18.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>122 </input>
<input>
<ID>IN_2</ID>114 </input>
<input>
<ID>IN_3</ID>106 </input>
<output>
<ID>OUT</ID>149 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-29.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT</ID>150 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-39</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>108 </input>
<output>
<ID>OUT</ID>151 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-50</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>117 </input>
<input>
<ID>IN_3</ID>109 </input>
<output>
<ID>OUT</ID>152 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-61</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT</ID>153 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-71.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>119 </input>
<input>
<ID>IN_3</ID>111 </input>
<output>
<ID>OUT</ID>154 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-82.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>112 </input>
<output>
<ID>OUT</ID>155 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>103</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>167,-51</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>151 </input>
<input>
<ID>IN_5</ID>150 </input>
<input>
<ID>IN_6</ID>149 </input>
<input>
<ID>IN_7</ID>148 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>75,-29.5</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>DD_KEYPAD_HEX</type>
<position>92.5,-36</position>
<output>
<ID>OUT_0</ID>161 </output>
<output>
<ID>OUT_1</ID>160 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>158 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>106</ID>
<type>DD_KEYPAD_HEX</type>
<position>92.5,-48</position>
<output>
<ID>OUT_0</ID>165 </output>
<output>
<ID>OUT_1</ID>164 </output>
<output>
<ID>OUT_2</ID>163 </output>
<output>
<ID>OUT_3</ID>162 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>92.5,-29</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>BA_DECODER_2x4</type>
<position>94.5,-3</position>
<input>
<ID>ENABLE</ID>170 </input>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT_0</ID>166 </output>
<output>
<ID>OUT_1</ID>167 </output>
<output>
<ID>OUT_2</ID>168 </output>
<output>
<ID>OUT_3</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>88.5,-2.5</position>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>86,-1</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>DD_KEYPAD_HEX</type>
<position>89.5,-15.5</position>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>172 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>90,-8.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AE_REGISTER8</type>
<position>109.5,-18.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>110 </output>
<output>
<ID>OUT_3</ID>109 </output>
<output>
<ID>OUT_4</ID>108 </output>
<output>
<ID>OUT_5</ID>107 </output>
<output>
<ID>OUT_6</ID>106 </output>
<output>
<ID>OUT_7</ID>105 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>166 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_REGISTER8</type>
<position>109.5,-31.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>120 </output>
<output>
<ID>OUT_1</ID>119 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>117 </output>
<output>
<ID>OUT_4</ID>116 </output>
<output>
<ID>OUT_5</ID>115 </output>
<output>
<ID>OUT_6</ID>114 </output>
<output>
<ID>OUT_7</ID>113 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>167 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>120,6</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-108,66,-100</points>
<connection>
<GID>9</GID>
<name>ENABLE_0</name></connection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-100,66,-100</points>
<connection>
<GID>1</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-98,64.5,-91.5</points>
<connection>
<GID>1</GID>
<name>write_clock</name></connection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-91.5,64.5,-91.5</points>
<connection>
<GID>16</GID>
<name>CLK</name></connection>
<intersection>28 11</intersection>
<intersection>64.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>28,-107,28,-91.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-91.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-116.5,63,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_0</name></connection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-116.5,64,-116.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-115.5,62,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_1</name></connection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-115.5,64,-115.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-114.5,61,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_2</name></connection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-114.5,64,-114.5</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-113.5,60,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_3</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-113.5,64,-113.5</points>
<connection>
<GID>9</GID>
<name>IN_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-112.5,59,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_4</name></connection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-112.5,64,-112.5</points>
<connection>
<GID>9</GID>
<name>IN_4</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-111.5,58,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_5</name></connection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-111.5,64,-111.5</points>
<connection>
<GID>9</GID>
<name>IN_5</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-110.5,57,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_6</name></connection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-110.5,64,-110.5</points>
<connection>
<GID>9</GID>
<name>IN_6</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-109.5,56,-106.5</points>
<connection>
<GID>1</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>1</GID>
<name>DATA_IN_7</name></connection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-109.5,64,-109.5</points>
<connection>
<GID>9</GID>
<name>IN_7</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-116.5,68.5,-115</points>
<intersection>-116.5 2</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-115,83.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>83.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-116.5,68.5,-116.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83.5,-115,83.5,-113</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115.5,68.5,-115</points>
<intersection>-115.5 2</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-115,81.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>81.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-115.5,68.5,-115.5</points>
<connection>
<GID>9</GID>
<name>OUT_1</name></connection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81.5,-115,81.5,-113</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115,68.5,-114.5</points>
<intersection>-115 1</intersection>
<intersection>-114.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-115,79.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>79.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-114.5,68.5,-114.5</points>
<connection>
<GID>9</GID>
<name>OUT_2</name></connection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>79.5,-115,79.5,-113</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-115,77.5,-115</points>
<intersection>68.5 3</intersection>
<intersection>77.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68.5,-115,68.5,-113.5</points>
<intersection>-115 1</intersection>
<intersection>-113.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>77.5,-115,77.5,-113</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>68,-113.5,68.5,-113.5</points>
<connection>
<GID>9</GID>
<name>OUT_3</name></connection>
<intersection>68.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115,68.5,-112.5</points>
<intersection>-115 1</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-115,75.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>75.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-112.5,68.5,-112.5</points>
<connection>
<GID>9</GID>
<name>OUT_4</name></connection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-115,75.5,-113</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115,68.5,-111.5</points>
<intersection>-115 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-111.5,68.5,-111.5</points>
<connection>
<GID>9</GID>
<name>OUT_5</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-115,73.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>73.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,-115,73.5,-113</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>-115 2</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115,68.5,-110.5</points>
<intersection>-115 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-115,71.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>71.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-110.5,68.5,-110.5</points>
<connection>
<GID>9</GID>
<name>OUT_6</name></connection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,-115,71.5,-113</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>-115 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-115,68.5,-109.5</points>
<intersection>-115 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-109.5,68.5,-109.5</points>
<connection>
<GID>9</GID>
<name>OUT_7</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-115,69.5,-115</points>
<intersection>68.5 0</intersection>
<intersection>69.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69.5,-115,69.5,-113</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<intersection>-115 2</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-96,54.5,-96</points>
<connection>
<GID>55</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-101,54.5,-101</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-103,54.5,-103</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-99,54.5,-99</points>
<connection>
<GID>55</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-100,54.5,-100</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-98,54.5,-98</points>
<connection>
<GID>55</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-102,54.5,-102</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-97,54.5,-97</points>
<connection>
<GID>55</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-108,40,-105</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-108,40,-108</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-14.5,131.5,-14.5</points>
<connection>
<GID>113</GID>
<name>OUT_7</name></connection>
<intersection>131.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131.5,-14.5,131.5,-4.5</points>
<intersection>-14.5 1</intersection>
<intersection>-4.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>131.5,-4.5,144.5,-4.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<intersection>131.5 4</intersection>
<intersection>143 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>143,-10.5,143,-4.5</points>
<intersection>-10.5 8</intersection>
<intersection>-4.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>143,-10.5,144.5,-10.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>143 6</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-15.5,144.5,-15.5</points>
<connection>
<GID>113</GID>
<name>OUT_6</name></connection>
<connection>
<GID>93</GID>
<name>IN_3</name></connection>
<connection>
<GID>61</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-26.5,130.5,-16.5</points>
<intersection>-26.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-26.5,144.5,-26.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<connection>
<GID>94</GID>
<name>IN_3</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-16.5,130.5,-16.5</points>
<connection>
<GID>113</GID>
<name>OUT_5</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-36,130,-17.5</points>
<intersection>-36 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-36,144.5,-36</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<connection>
<GID>98</GID>
<name>IN_3</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-17.5,130,-17.5</points>
<connection>
<GID>113</GID>
<name>OUT_4</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-47,129.5,-18.5</points>
<intersection>-47 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-47,144.5,-47</points>
<connection>
<GID>64</GID>
<name>IN_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_3</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-18.5,129.5,-18.5</points>
<connection>
<GID>113</GID>
<name>OUT_3</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-58,129,-19.5</points>
<intersection>-58 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-58,144.5,-58</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-19.5,129,-19.5</points>
<connection>
<GID>113</GID>
<name>OUT_2</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-68.5,128.5,-20.5</points>
<intersection>-68.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-68.5,144.5,-68.5</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-20.5,128.5,-20.5</points>
<connection>
<GID>113</GID>
<name>OUT_1</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-79.5,128,-21.5</points>
<intersection>-79.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-21.5,128,-21.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-79.5,144.5,-79.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-27.5,127,-6.5</points>
<intersection>-27.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-6.5,144.5,-6.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-27.5,127,-27.5</points>
<connection>
<GID>114</GID>
<name>OUT_7</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-28.5,126.5,-17.5</points>
<intersection>-28.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-17.5,144.5,-17.5</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<connection>
<GID>93</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-28.5,126.5,-28.5</points>
<connection>
<GID>114</GID>
<name>OUT_6</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-29.5,132,-29.5</points>
<connection>
<GID>114</GID>
<name>OUT_5</name></connection>
<intersection>132 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132,-29.5,132,-28.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-29.5 1</intersection>
<intersection>-28.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>132,-28.5,144.5,-28.5</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>132 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-38,126,-30.5</points>
<intersection>-38 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-38,144.5,-38</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-30.5,126,-30.5</points>
<connection>
<GID>114</GID>
<name>OUT_4</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-49,125.5,-31.5</points>
<intersection>-49 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-49,144.5,-49</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-31.5,125.5,-31.5</points>
<connection>
<GID>114</GID>
<name>OUT_3</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-60,125,-32.5</points>
<intersection>-60 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-60,144.5,-60</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-32.5,125,-32.5</points>
<connection>
<GID>114</GID>
<name>OUT_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-70.5,124.5,-33.5</points>
<intersection>-70.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-33.5,124.5,-33.5</points>
<connection>
<GID>114</GID>
<name>OUT_1</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-70.5,144.5,-70.5</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-81.5,127.5,-34.5</points>
<intersection>-81.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-81.5,144.5,-81.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-34.5,127.5,-34.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-41,123,-8.5</points>
<intersection>-41 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-8.5,144.5,-8.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-41,123,-41</points>
<connection>
<GID>58</GID>
<name>OUT_7</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-42,122.5,-19.5</points>
<intersection>-42 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-19.5,144.5,-19.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-42,122.5,-42</points>
<connection>
<GID>58</GID>
<name>OUT_6</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-43,122,-30.5</points>
<intersection>-43 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-30.5,144.5,-30.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-43,122,-43</points>
<connection>
<GID>58</GID>
<name>OUT_5</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-44,121.5,-40</points>
<intersection>-44 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-40,144.5,-40</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-44,121.5,-44</points>
<connection>
<GID>58</GID>
<name>OUT_4</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-51,121,-45</points>
<intersection>-51 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-51,144.5,-51</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-45,121,-45</points>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-62,120.5,-46</points>
<intersection>-62 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-62,144.5,-62</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-46,120.5,-46</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-72.5,120,-47</points>
<intersection>-72.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-72.5,144.5,-72.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-47,120,-47</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-83.5,119.5,-48</points>
<intersection>-83.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-48,119.5,-48</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-83.5,144.5,-83.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-54,118.5,-10.5</points>
<intersection>-54 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-10.5,132,-10.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-54,118.5,-54</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-55,118,-21.5</points>
<intersection>-55 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-21.5,144.5,-21.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-55,118,-55</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-56,117.5,-32.5</points>
<intersection>-56 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-32.5,144.5,-32.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-56,117.5,-56</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-42,144.5,-42</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113.5,-57,113.5,-42</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-58,116.5,-53</points>
<intersection>-58 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-53,144.5,-53</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-58,116.5,-58</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-64,116,-59</points>
<intersection>-64 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-64,144.5,-64</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-59,116,-59</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-74.5,115.5,-60</points>
<intersection>-74.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-74.5,144.5,-74.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-60,115.5,-60</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-36,156.5,-7.5</points>
<intersection>-36 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-7.5,156.5,-7.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-36,162,-36</points>
<connection>
<GID>70</GID>
<name>IN_7</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-37,156.5,-18.5</points>
<intersection>-37 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-18.5,156.5,-18.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-37,162,-37</points>
<connection>
<GID>70</GID>
<name>IN_6</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-38,156.5,-29.5</points>
<intersection>-38 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-29.5,156.5,-29.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-38,162,-38</points>
<connection>
<GID>70</GID>
<name>IN_5</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,-39,162,-39</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-50,156.5,-40</points>
<intersection>-50 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-50,156.5,-50</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-40,162,-40</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-61,156.5,-41</points>
<intersection>-61 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-61,156.5,-61</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-41,162,-41</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-71.5,156.5,-42</points>
<intersection>-71.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-71.5,156.5,-71.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-42,162,-42</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-82.5,156.5,-43</points>
<intersection>-82.5 2</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-43,162,-43</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-82.5,156.5,-82.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-85.5,115,-61</points>
<intersection>-85.5 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-85.5,144.5,-85.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-61,115,-61</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-66.5,105,-23.5</points>
<intersection>-66.5 10</intersection>
<intersection>-63 8</intersection>
<intersection>-50 7</intersection>
<intersection>-36.5 6</intersection>
<intersection>-23.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>105,-23.5,108.5,-23.5</points>
<connection>
<GID>113</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105,-36.5,108.5,-36.5</points>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>105,-50,108.5,-50</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>105,-63,108.5,-63</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-66.5,105,-66.5</points>
<connection>
<GID>72</GID>
<name>CLK</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-77.5,136,0.5</points>
<connection>
<GID>69</GID>
<name>SEL_0</name></connection>
<connection>
<GID>66</GID>
<name>SEL_0</name></connection>
<connection>
<GID>65</GID>
<name>SEL_0</name></connection>
<connection>
<GID>64</GID>
<name>SEL_0</name></connection>
<connection>
<GID>63</GID>
<name>SEL_0</name></connection>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<connection>
<GID>61</GID>
<name>SEL_0</name></connection>
<connection>
<GID>60</GID>
<name>SEL_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,0.5,136,0.5</points>
<intersection>82.5 2</intersection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>82.5,-25.5,82.5,0.5</points>
<intersection>-25.5 3</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-25.5,82.5,-25.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>82.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-77.5,135,0</points>
<connection>
<GID>69</GID>
<name>SEL_1</name></connection>
<connection>
<GID>66</GID>
<name>SEL_1</name></connection>
<connection>
<GID>65</GID>
<name>SEL_1</name></connection>
<connection>
<GID>64</GID>
<name>SEL_1</name></connection>
<connection>
<GID>63</GID>
<name>SEL_1</name></connection>
<connection>
<GID>62</GID>
<name>SEL_1</name></connection>
<connection>
<GID>61</GID>
<name>SEL_1</name></connection>
<connection>
<GID>60</GID>
<name>SEL_1</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,0,135,0</points>
<intersection>82 2</intersection>
<intersection>135 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>82,-23.5,82,0</points>
<intersection>-23.5 3</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-23.5,82,-23.5</points>
<connection>
<GID>71</GID>
<name>OUT_1</name></connection>
<intersection>82 2</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-47,151,-7.5</points>
<intersection>-47 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-7.5,151,-7.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-47,162,-47</points>
<connection>
<GID>103</GID>
<name>IN_7</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-48,151,-18.5</points>
<intersection>-48 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-18.5,151,-18.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-48,162,-48</points>
<connection>
<GID>103</GID>
<name>IN_6</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-49,151,-29.5</points>
<intersection>-49 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-29.5,151,-29.5</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-49,162,-49</points>
<connection>
<GID>103</GID>
<name>IN_5</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-50,151,-39</points>
<intersection>-50 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-39,151,-39</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-50,162,-50</points>
<connection>
<GID>103</GID>
<name>IN_4</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-51,162,-51</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-51,151,-50</points>
<intersection>-51 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150.5,-50,151,-50</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-61,151,-52</points>
<intersection>-61 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-61,151,-61</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-52,162,-52</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-71.5,151,-53</points>
<intersection>-71.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-71.5,151,-71.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-53,162,-53</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-82.5,151,-54</points>
<intersection>-82.5 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-54,162,-54</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150.5,-82.5,151,-82.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-77.5,148.5,-1</points>
<connection>
<GID>102</GID>
<name>SEL_0</name></connection>
<connection>
<GID>101</GID>
<name>SEL_0</name></connection>
<connection>
<GID>100</GID>
<name>SEL_0</name></connection>
<connection>
<GID>99</GID>
<name>SEL_0</name></connection>
<connection>
<GID>98</GID>
<name>SEL_0</name></connection>
<connection>
<GID>94</GID>
<name>SEL_0</name></connection>
<connection>
<GID>93</GID>
<name>SEL_0</name></connection>
<connection>
<GID>87</GID>
<name>SEL_0</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-1,148.5,-1</points>
<intersection>83.5 2</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,-39.5,83.5,-1</points>
<intersection>-39.5 3</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-39.5,83.5,-39.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>83.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-77.5,147.5,-0.5</points>
<connection>
<GID>102</GID>
<name>SEL_1</name></connection>
<connection>
<GID>101</GID>
<name>SEL_1</name></connection>
<connection>
<GID>100</GID>
<name>SEL_1</name></connection>
<connection>
<GID>99</GID>
<name>SEL_1</name></connection>
<connection>
<GID>98</GID>
<name>SEL_1</name></connection>
<connection>
<GID>94</GID>
<name>SEL_1</name></connection>
<connection>
<GID>93</GID>
<name>SEL_1</name></connection>
<connection>
<GID>87</GID>
<name>SEL_1</name></connection>
<intersection>-0.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>83,-0.5,147.5,-0.5</points>
<intersection>83 16</intersection>
<intersection>147.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>83,-37.5,83,-0.5</points>
<intersection>-37.5 18</intersection>
<intersection>-0.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>81.5,-37.5,83,-37.5</points>
<connection>
<GID>78</GID>
<name>OUT_1</name></connection>
<intersection>83 16</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-54,104,-14.5</points>
<intersection>-54 6</intersection>
<intersection>-41 3</intersection>
<intersection>-33 4</intersection>
<intersection>-27.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-14.5,105.5,-14.5</points>
<connection>
<GID>113</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-27.5,105.5,-27.5</points>
<connection>
<GID>114</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-41,105.5,-41</points>
<connection>
<GID>58</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>97.5,-33,104,-33</points>
<connection>
<GID>105</GID>
<name>OUT_3</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104,-54,105.5,-54</points>
<connection>
<GID>59</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-55,103.5,-15.5</points>
<intersection>-55 6</intersection>
<intersection>-42 5</intersection>
<intersection>-35 2</intersection>
<intersection>-28.5 3</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-35,103.5,-35</points>
<connection>
<GID>105</GID>
<name>OUT_2</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-28.5,105.5,-28.5</points>
<connection>
<GID>114</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103.5,-15.5,105.5,-15.5</points>
<connection>
<GID>113</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103.5,-42,105.5,-42</points>
<connection>
<GID>58</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103.5,-55,105.5,-55</points>
<connection>
<GID>59</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-56,103,-16.5</points>
<intersection>-56 6</intersection>
<intersection>-43 3</intersection>
<intersection>-37 2</intersection>
<intersection>-29.5 4</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-37,103,-37</points>
<connection>
<GID>105</GID>
<name>OUT_1</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-43,105.5,-43</points>
<connection>
<GID>58</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103,-29.5,105.5,-29.5</points>
<connection>
<GID>114</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,-16.5,105.5,-16.5</points>
<connection>
<GID>113</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103,-56,105.5,-56</points>
<connection>
<GID>59</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-57,102.5,-17.5</points>
<intersection>-57 6</intersection>
<intersection>-44 3</intersection>
<intersection>-39 2</intersection>
<intersection>-30.5 4</intersection>
<intersection>-17.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-39,102.5,-39</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-44,105.5,-44</points>
<connection>
<GID>58</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102.5,-30.5,105.5,-30.5</points>
<connection>
<GID>114</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102.5,-17.5,105.5,-17.5</points>
<connection>
<GID>113</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102.5,-57,105.5,-57</points>
<connection>
<GID>59</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-58,102,-18.5</points>
<intersection>-58 5</intersection>
<intersection>-45 2</intersection>
<intersection>-31.5 3</intersection>
<intersection>-18.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-45,105.5,-45</points>
<connection>
<GID>58</GID>
<name>IN_3</name></connection>
<connection>
<GID>106</GID>
<name>OUT_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-31.5,105.5,-31.5</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102,-18.5,105.5,-18.5</points>
<connection>
<GID>113</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102,-58,105.5,-58</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-59,101.5,-19.5</points>
<intersection>-59 5</intersection>
<intersection>-47 2</intersection>
<intersection>-46 4</intersection>
<intersection>-32.5 3</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-19.5,105.5,-19.5</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-47,101.5,-47</points>
<connection>
<GID>106</GID>
<name>OUT_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-32.5,105.5,-32.5</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101.5,-46,105.5,-46</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101.5,-59,105.5,-59</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-60,101,-20.5</points>
<intersection>-60 5</intersection>
<intersection>-49 2</intersection>
<intersection>-47 4</intersection>
<intersection>-33.5 3</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-20.5,105.5,-20.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-49,101,-49</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-33.5,105.5,-33.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101,-47,105.5,-47</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101,-60,105.5,-60</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-61,100.5,-21.5</points>
<intersection>-61 5</intersection>
<intersection>-51 2</intersection>
<intersection>-48 4</intersection>
<intersection>-34.5 3</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-21.5,105.5,-21.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-51,100.5,-51</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-34.5,105.5,-34.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>100.5,-48,105.5,-48</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>100.5,-61,105.5,-61</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-12.5,107.5,-4.5</points>
<intersection>-12.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-4.5,107.5,-4.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-12.5,108.5,-12.5</points>
<connection>
<GID>113</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-25.5,107.5,-3.5</points>
<intersection>-25.5 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-3.5,107.5,-3.5</points>
<connection>
<GID>108</GID>
<name>OUT_1</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-25.5,108.5,-25.5</points>
<connection>
<GID>114</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-39,107.5,-2.5</points>
<intersection>-39 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-2.5,107.5,-2.5</points>
<connection>
<GID>108</GID>
<name>OUT_2</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-39,108.5,-39</points>
<connection>
<GID>58</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-52,107.5,-1.5</points>
<intersection>-52 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-1.5,107.5,-1.5</points>
<connection>
<GID>108</GID>
<name>OUT_3</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-52,108.5,-52</points>
<connection>
<GID>59</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-2.5,91.5,-2.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>91.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91.5,-2.5,91.5,-1.5</points>
<connection>
<GID>108</GID>
<name>ENABLE</name></connection>
<intersection>-2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-18.5,96,-7.5</points>
<intersection>-18.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-7.5,96,-7.5</points>
<intersection>91 3</intersection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-18.5,96,-18.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91,-7.5,91,-4.5</points>
<intersection>-7.5 1</intersection>
<intersection>-4.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>91,-4.5,91.5,-4.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>91 3</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-16.5,96.5,-7</points>
<intersection>-16.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-7,96.5,-7</points>
<intersection>91.5 3</intersection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-16.5,96.5,-16.5</points>
<connection>
<GID>111</GID>
<name>OUT_1</name></connection>
<intersection>96.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-7,91.5,-3.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>63.675,150.224,1841.68,-766.776</PageViewport>
<gate>
<ID>196</ID>
<type>AA_INVERTER</type>
<position>70,-67.5</position>
<input>
<ID>IN_0</ID>268 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>94.5,-43</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>72,-75</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>72,-76.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AE_REGISTER8</type>
<position>99,-59</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>174 </input>
<input>
<ID>IN_2</ID>175 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_4</ID>177 </input>
<input>
<ID>IN_5</ID>178 </input>
<input>
<ID>IN_6</ID>179 </input>
<input>
<ID>IN_7</ID>180 </input>
<output>
<ID>OUT_0</ID>188 </output>
<output>
<ID>OUT_1</ID>187 </output>
<output>
<ID>OUT_2</ID>186 </output>
<output>
<ID>OUT_3</ID>185 </output>
<output>
<ID>OUT_4</ID>184 </output>
<output>
<ID>OUT_5</ID>183 </output>
<output>
<ID>OUT_6</ID>182 </output>
<output>
<ID>OUT_7</ID>181 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>267 </input>
<input>
<ID>count_enable</ID>203 </input>
<input>
<ID>count_up</ID>203 </input>
<input>
<ID>load</ID>269 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_REGISTER8</type>
<position>116,-59</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>186 </input>
<input>
<ID>IN_3</ID>185 </input>
<input>
<ID>IN_4</ID>184 </input>
<input>
<ID>IN_5</ID>183 </input>
<input>
<ID>IN_6</ID>182 </input>
<input>
<ID>IN_7</ID>181 </input>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>217 </output>
<output>
<ID>OUT_2</ID>194 </output>
<output>
<ID>OUT_3</ID>193 </output>
<output>
<ID>OUT_4</ID>192 </output>
<output>
<ID>OUT_5</ID>191 </output>
<output>
<ID>OUT_6</ID>190 </output>
<output>
<ID>OUT_7</ID>189 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>202 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_REGISTER8</type>
<position>153,-76.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>256 </input>
<input>
<ID>IN_2</ID>257 </input>
<input>
<ID>IN_3</ID>258 </input>
<input>
<ID>IN_4</ID>259 </input>
<input>
<ID>IN_5</ID>254 </input>
<input>
<ID>IN_6</ID>261 </input>
<input>
<ID>IN_7</ID>260 </input>
<output>
<ID>OUT_0</ID>226 </output>
<output>
<ID>OUT_1</ID>225 </output>
<output>
<ID>OUT_2</ID>224 </output>
<output>
<ID>OUT_3</ID>223 </output>
<output>
<ID>OUT_4</ID>222 </output>
<output>
<ID>OUT_5</ID>221 </output>
<output>
<ID>OUT_6</ID>220 </output>
<output>
<ID>OUT_7</ID>219 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>216 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_RAM_8x8</type>
<position>131,-58.5</position>
<input>
<ID>ADDRESS_0</ID>218 </input>
<input>
<ID>ADDRESS_1</ID>217 </input>
<input>
<ID>ADDRESS_2</ID>194 </input>
<input>
<ID>ADDRESS_3</ID>193 </input>
<input>
<ID>ADDRESS_4</ID>192 </input>
<input>
<ID>ADDRESS_5</ID>191 </input>
<input>
<ID>ADDRESS_6</ID>190 </input>
<input>
<ID>ADDRESS_7</ID>189 </input>
<input>
<ID>DATA_IN_0</ID>262 </input>
<input>
<ID>DATA_IN_1</ID>242 </input>
<input>
<ID>DATA_IN_2</ID>245 </input>
<input>
<ID>DATA_IN_3</ID>246 </input>
<input>
<ID>DATA_IN_4</ID>247 </input>
<input>
<ID>DATA_IN_5</ID>251 </input>
<input>
<ID>DATA_IN_6</ID>252 </input>
<input>
<ID>DATA_IN_7</ID>253 </input>
<output>
<ID>DATA_OUT_0</ID>262 </output>
<output>
<ID>DATA_OUT_1</ID>242 </output>
<output>
<ID>DATA_OUT_2</ID>245 </output>
<output>
<ID>DATA_OUT_3</ID>246 </output>
<output>
<ID>DATA_OUT_4</ID>247 </output>
<output>
<ID>DATA_OUT_5</ID>251 </output>
<output>
<ID>DATA_OUT_6</ID>252 </output>
<output>
<ID>DATA_OUT_7</ID>253 </output>
<input>
<ID>ENABLE_0</ID>241 </input>
<input>
<ID>write_enable</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 170</lparam>
<lparam>Address:1 187</lparam>
<lparam>Address:2 204</lparam>
<lparam>Address:3 221</lparam></gate>
<gate>
<ID>127</ID>
<type>AE_REGISTER8</type>
<position>169,-76.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>225 </input>
<input>
<ID>IN_2</ID>224 </input>
<input>
<ID>IN_3</ID>223 </input>
<input>
<ID>IN_4</ID>222 </input>
<input>
<ID>IN_5</ID>221 </input>
<input>
<ID>IN_6</ID>220 </input>
<input>
<ID>IN_7</ID>219 </input>
<output>
<ID>OUT_0</ID>236 </output>
<output>
<ID>OUT_1</ID>237 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>227 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>131</ID>
<type>DD_KEYPAD_HEX</type>
<position>79.5,-65</position>
<output>
<ID>OUT_0</ID>173 </output>
<output>
<ID>OUT_1</ID>174 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>176 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>133</ID>
<type>DD_KEYPAD_HEX</type>
<position>79.5,-53</position>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>178 </output>
<output>
<ID>OUT_2</ID>179 </output>
<output>
<ID>OUT_3</ID>180 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>135</ID>
<type>BB_CLOCK</type>
<position>68,-90.5</position>
<output>
<ID>CLK</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>97,-40</position>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>84.5,-42</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>84.5,-39.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>110,-42.5</position>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>98,-87.5</position>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>92.5,-84.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>149,-69</position>
<output>
<ID>OUT_0</ID>216 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>94,-51</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>110.5,-51</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>131,-50</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>153,-66</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>166,-68.5</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>169</ID>
<type>BE_ROM_8x8</type>
<position>184,-76</position>
<input>
<ID>ADDRESS_0</ID>236 </input>
<input>
<ID>ADDRESS_1</ID>237 </input>
<input>
<ID>ENABLE_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>141,-56</position>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>141,-59</position>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>147.5,-55.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>148,-58.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>145,-76</position>
<input>
<ID>ENABLE_0</ID>241 </input>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>245 </input>
<input>
<ID>IN_3</ID>246 </input>
<input>
<ID>IN_4</ID>247 </input>
<input>
<ID>IN_5</ID>251 </input>
<input>
<ID>IN_6</ID>252 </input>
<input>
<ID>IN_7</ID>253 </input>
<output>
<ID>OUT_0</ID>255 </output>
<output>
<ID>OUT_1</ID>256 </output>
<output>
<ID>OUT_2</ID>257 </output>
<output>
<ID>OUT_3</ID>258 </output>
<output>
<ID>OUT_4</ID>259 </output>
<output>
<ID>OUT_5</ID>254 </output>
<output>
<ID>OUT_6</ID>261 </output>
<output>
<ID>OUT_7</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>178</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>124,-76</position>
<input>
<ID>ENABLE_0</ID>240 </input>
<output>
<ID>OUT_0</ID>262 </output>
<output>
<ID>OUT_1</ID>242 </output>
<output>
<ID>OUT_2</ID>245 </output>
<output>
<ID>OUT_3</ID>246 </output>
<output>
<ID>OUT_4</ID>247 </output>
<output>
<ID>OUT_5</ID>251 </output>
<output>
<ID>OUT_6</ID>252 </output>
<output>
<ID>OUT_7</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>170.5,-68</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>193,-76.5</position>
<output>
<ID>OUT_0</ID>264 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>194.5,-73.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_AND2</type>
<position>94,-72</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>79.5,-89.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>74,-86.5</position>
<output>
<ID>OUT_0</ID>266 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>65,-73</position>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-59,126,-59</points>
<connection>
<GID>119</GID>
<name>OUT_3</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-60,126,-60</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-53,115,-42.5</points>
<connection>
<GID>119</GID>
<name>load</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-42.5,115,-42.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-53,99,-40</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>count_enable</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99,-52,100,-52</points>
<intersection>99 0</intersection>
<intersection>100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100,-53,100,-52</points>
<connection>
<GID>117</GID>
<name>count_up</name></connection>
<intersection>-52 2</intersection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>151,-69,152,-69</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>152 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>152,-70.5,152,-69</points>
<connection>
<GID>123</GID>
<name>load</name></connection>
<intersection>-69 2</intersection></vsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-61,126,-61</points>
<connection>
<GID>119</GID>
<name>OUT_1</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-62,126,-62</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-72.5,165,-72.5</points>
<connection>
<GID>123</GID>
<name>OUT_7</name></connection>
<connection>
<GID>127</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-73.5,165,-73.5</points>
<connection>
<GID>123</GID>
<name>OUT_6</name></connection>
<connection>
<GID>127</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-74.5,165,-74.5</points>
<connection>
<GID>123</GID>
<name>OUT_5</name></connection>
<connection>
<GID>127</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-75.5,165,-75.5</points>
<connection>
<GID>123</GID>
<name>OUT_4</name></connection>
<connection>
<GID>127</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-76.5,165,-76.5</points>
<connection>
<GID>123</GID>
<name>OUT_3</name></connection>
<connection>
<GID>127</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-77.5,165,-77.5</points>
<connection>
<GID>123</GID>
<name>OUT_2</name></connection>
<connection>
<GID>127</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-78.5,165,-78.5</points>
<connection>
<GID>123</GID>
<name>OUT_1</name></connection>
<connection>
<GID>127</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-79.5,165,-79.5</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-70.5,168,-68.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173,-79.5,179,-79.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<connection>
<GID>169</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173,-78.5,179,-78.5</points>
<connection>
<GID>127</GID>
<name>OUT_1</name></connection>
<connection>
<GID>169</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-89.5,115,-64</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-89.5,168,-89.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>85 6</intersection>
<intersection>115 0</intersection>
<intersection>152 5</intersection>
<intersection>168 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>168,-89.5,168,-81.5</points>
<connection>
<GID>127</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>152,-89.5,152,-81.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>85,-89.5,85,-71</points>
<intersection>-89.5 1</intersection>
<intersection>-71 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>85,-71,91,-71</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>85 6</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-87.5,100,-64</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,-87.5,170,-87.5</points>
<intersection>100 0</intersection>
<intersection>117 3</intersection>
<intersection>154 7</intersection>
<intersection>170 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-87.5,117,-64</points>
<connection>
<GID>119</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>170,-87.5,170,-81.5</points>
<connection>
<GID>127</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>154,-87.5,154,-81.5</points>
<connection>
<GID>123</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-56,139,-56</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>136 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>136,-71,136,-56</points>
<connection>
<GID>125</GID>
<name>write_enable</name></connection>
<intersection>-71 4</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,-71,136,-71</points>
<connection>
<GID>178</GID>
<name>ENABLE_0</name></connection>
<intersection>136 3</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-59,139,-59</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ENABLE_0</name></connection>
<intersection>139 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>139,-71,139,-59</points>
<intersection>-71 6</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-71,145,-71</points>
<connection>
<GID>177</GID>
<name>ENABLE_0</name></connection>
<intersection>139 5</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-78.5,143,-78.5</points>
<connection>
<GID>178</GID>
<name>OUT_1</name></connection>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>133.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>133.5,-78.5,133.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-77.5,143,-77.5</points>
<connection>
<GID>178</GID>
<name>OUT_2</name></connection>
<connection>
<GID>177</GID>
<name>IN_2</name></connection>
<intersection>132.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132.5,-77.5,132.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_2</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-76.5,143,-76.5</points>
<connection>
<GID>178</GID>
<name>OUT_3</name></connection>
<connection>
<GID>177</GID>
<name>IN_3</name></connection>
<intersection>131.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>131.5,-76.5,131.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_3</name></connection>
<intersection>-76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-75.5,143,-75.5</points>
<connection>
<GID>178</GID>
<name>OUT_4</name></connection>
<connection>
<GID>177</GID>
<name>IN_4</name></connection>
<intersection>130.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130.5,-75.5,130.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_4</name></connection>
<intersection>-75.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-74.5,143,-74.5</points>
<connection>
<GID>178</GID>
<name>OUT_5</name></connection>
<connection>
<GID>177</GID>
<name>IN_5</name></connection>
<intersection>129.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>129.5,-74.5,129.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_5</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-73.5,143,-73.5</points>
<connection>
<GID>178</GID>
<name>OUT_6</name></connection>
<connection>
<GID>177</GID>
<name>IN_6</name></connection>
<intersection>128.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-73.5,128.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_6</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-72.5,143,-72.5</points>
<connection>
<GID>178</GID>
<name>OUT_7</name></connection>
<connection>
<GID>177</GID>
<name>IN_7</name></connection>
<intersection>127.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127.5,-72.5,127.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_7</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-74.5,149,-74.5</points>
<connection>
<GID>123</GID>
<name>IN_5</name></connection>
<connection>
<GID>177</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-79.5,149,-79.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-78.5,149,-78.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<connection>
<GID>177</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-77.5,149,-77.5</points>
<connection>
<GID>123</GID>
<name>IN_2</name></connection>
<connection>
<GID>177</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-76.5,149,-76.5</points>
<connection>
<GID>123</GID>
<name>IN_3</name></connection>
<connection>
<GID>177</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-75.5,149,-75.5</points>
<connection>
<GID>123</GID>
<name>IN_4</name></connection>
<connection>
<GID>177</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-72.5,149,-72.5</points>
<connection>
<GID>123</GID>
<name>IN_7</name></connection>
<connection>
<GID>177</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-73.5,149,-73.5</points>
<connection>
<GID>123</GID>
<name>IN_6</name></connection>
<connection>
<GID>177</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-79.5,143,-79.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>134.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-79.5,134.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_0</name></connection>
<intersection>-79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-76.5,191,-76.5</points>
<connection>
<GID>169</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-90.5,76.5,-90.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-88.5,76.5,-86.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-86.5,76.5,-86.5</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-72,98,-64</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-72,98,-72</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-73,91,-73</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>70 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>70,-73,70,-70.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-53,98,-45</points>
<connection>
<GID>117</GID>
<name>load</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-64.5,70,-45</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-45,98,-45</points>
<intersection>70 1</intersection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-68,89.5,-62</points>
<intersection>-68 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-62,95,-62</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-68,89.5,-68</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-66,89.5,-61</points>
<intersection>-66 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-61,95,-61</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-66,89.5,-66</points>
<connection>
<GID>131</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-64,89.5,-60</points>
<intersection>-64 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-60,95,-60</points>
<connection>
<GID>117</GID>
<name>IN_2</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-64,89.5,-64</points>
<connection>
<GID>131</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-62,89.5,-59</points>
<intersection>-62 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-59,95,-59</points>
<connection>
<GID>117</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-62,89.5,-62</points>
<connection>
<GID>131</GID>
<name>OUT_3</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-58,89.5,-56</points>
<intersection>-58 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-58,95,-58</points>
<connection>
<GID>117</GID>
<name>IN_4</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-56,89.5,-56</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-57,89.5,-54</points>
<intersection>-57 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-57,95,-57</points>
<connection>
<GID>117</GID>
<name>IN_5</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-54,89.5,-54</points>
<connection>
<GID>133</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-56,89.5,-52</points>
<intersection>-56 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-56,95,-56</points>
<connection>
<GID>117</GID>
<name>IN_6</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-52,89.5,-52</points>
<connection>
<GID>133</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-55,95,-55</points>
<connection>
<GID>117</GID>
<name>IN_7</name></connection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-55,84.5,-50</points>
<connection>
<GID>133</GID>
<name>OUT_3</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-55,112,-55</points>
<connection>
<GID>119</GID>
<name>IN_7</name></connection>
<connection>
<GID>117</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-56,112,-56</points>
<connection>
<GID>119</GID>
<name>IN_6</name></connection>
<connection>
<GID>117</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-57,112,-57</points>
<connection>
<GID>119</GID>
<name>IN_5</name></connection>
<connection>
<GID>117</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-58,112,-58</points>
<connection>
<GID>119</GID>
<name>IN_4</name></connection>
<connection>
<GID>117</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-59,112,-59</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<connection>
<GID>117</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-60,112,-60</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<connection>
<GID>117</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-61,112,-61</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>117</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-62,112,-62</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-55,126,-55</points>
<connection>
<GID>119</GID>
<name>OUT_7</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-56,126,-56</points>
<connection>
<GID>119</GID>
<name>OUT_6</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-57,126,-57</points>
<connection>
<GID>119</GID>
<name>OUT_5</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-58,126,-58</points>
<connection>
<GID>119</GID>
<name>OUT_4</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-70.0998,627.373,1707.9,-289.627</PageViewport>
<gate>
<ID>204</ID>
<type>AA_INVERTER</type>
<position>50.5,-52.5</position>
<input>
<ID>IN_0</ID>333 </input>
<output>
<ID>OUT_0</ID>334 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_TOGGLE</type>
<position>75,-28</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>52.5,-60</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>52.5,-61.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AE_REGISTER8</type>
<position>79.5,-44</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>272 </input>
<input>
<ID>IN_2</ID>273 </input>
<input>
<ID>IN_3</ID>274 </input>
<input>
<ID>IN_4</ID>275 </input>
<input>
<ID>IN_5</ID>276 </input>
<input>
<ID>IN_6</ID>277 </input>
<input>
<ID>IN_7</ID>278 </input>
<output>
<ID>OUT_0</ID>286 </output>
<output>
<ID>OUT_1</ID>285 </output>
<output>
<ID>OUT_2</ID>284 </output>
<output>
<ID>OUT_3</ID>283 </output>
<output>
<ID>OUT_4</ID>282 </output>
<output>
<ID>OUT_5</ID>281 </output>
<output>
<ID>OUT_6</ID>280 </output>
<output>
<ID>OUT_7</ID>279 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>332 </input>
<input>
<ID>count_enable</ID>294 </input>
<input>
<ID>count_up</ID>294 </input>
<input>
<ID>load</ID>334 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>209</ID>
<type>AE_REGISTER8</type>
<position>96.5,-44</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>285 </input>
<input>
<ID>IN_2</ID>284 </input>
<input>
<ID>IN_3</ID>283 </input>
<input>
<ID>IN_4</ID>282 </input>
<input>
<ID>IN_5</ID>281 </input>
<input>
<ID>IN_6</ID>280 </input>
<input>
<ID>IN_7</ID>279 </input>
<output>
<ID>OUT_0</ID>297 </output>
<output>
<ID>OUT_1</ID>296 </output>
<output>
<ID>OUT_2</ID>292 </output>
<output>
<ID>OUT_3</ID>291 </output>
<output>
<ID>OUT_4</ID>290 </output>
<output>
<ID>OUT_5</ID>289 </output>
<output>
<ID>OUT_6</ID>288 </output>
<output>
<ID>OUT_7</ID>287 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>309 </input>
<input>
<ID>load</ID>293 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_REGISTER8</type>
<position>133.5,-61.5</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>322 </input>
<input>
<ID>IN_2</ID>323 </input>
<input>
<ID>IN_3</ID>324 </input>
<input>
<ID>IN_4</ID>325 </input>
<input>
<ID>IN_5</ID>320 </input>
<input>
<ID>IN_6</ID>327 </input>
<input>
<ID>IN_7</ID>326 </input>
<output>
<ID>OUT_0</ID>305 </output>
<output>
<ID>OUT_1</ID>304 </output>
<output>
<ID>OUT_2</ID>303 </output>
<output>
<ID>OUT_3</ID>302 </output>
<output>
<ID>OUT_4</ID>301 </output>
<output>
<ID>OUT_5</ID>300 </output>
<output>
<ID>OUT_6</ID>299 </output>
<output>
<ID>OUT_7</ID>298 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>309 </input>
<input>
<ID>load</ID>295 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_RAM_8x8</type>
<position>111.5,-43.5</position>
<input>
<ID>ADDRESS_0</ID>297 </input>
<input>
<ID>ADDRESS_1</ID>296 </input>
<input>
<ID>ADDRESS_2</ID>292 </input>
<input>
<ID>ADDRESS_3</ID>291 </input>
<input>
<ID>ADDRESS_4</ID>290 </input>
<input>
<ID>ADDRESS_5</ID>289 </input>
<input>
<ID>ADDRESS_6</ID>288 </input>
<input>
<ID>ADDRESS_7</ID>287 </input>
<input>
<ID>DATA_IN_0</ID>328 </input>
<input>
<ID>DATA_IN_1</ID>313 </input>
<input>
<ID>DATA_IN_2</ID>314 </input>
<input>
<ID>DATA_IN_3</ID>315 </input>
<input>
<ID>DATA_IN_4</ID>316 </input>
<input>
<ID>DATA_IN_5</ID>317 </input>
<input>
<ID>DATA_IN_6</ID>318 </input>
<input>
<ID>DATA_IN_7</ID>319 </input>
<output>
<ID>DATA_OUT_0</ID>328 </output>
<output>
<ID>DATA_OUT_1</ID>313 </output>
<output>
<ID>DATA_OUT_2</ID>314 </output>
<output>
<ID>DATA_OUT_3</ID>315 </output>
<output>
<ID>DATA_OUT_4</ID>316 </output>
<output>
<ID>DATA_OUT_5</ID>317 </output>
<output>
<ID>DATA_OUT_6</ID>318 </output>
<output>
<ID>DATA_OUT_7</ID>319 </output>
<input>
<ID>ENABLE_0</ID>312 </input>
<input>
<ID>write_enable</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_REGISTER8</type>
<position>149.5,-61.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>304 </input>
<input>
<ID>IN_2</ID>303 </input>
<input>
<ID>IN_3</ID>302 </input>
<input>
<ID>IN_4</ID>301 </input>
<input>
<ID>IN_5</ID>300 </input>
<input>
<ID>IN_6</ID>299 </input>
<input>
<ID>IN_7</ID>298 </input>
<output>
<ID>OUT_0</ID>307 </output>
<output>
<ID>OUT_1</ID>308 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>309 </input>
<input>
<ID>load</ID>306 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>213</ID>
<type>DD_KEYPAD_HEX</type>
<position>60,-50</position>
<output>
<ID>OUT_0</ID>271 </output>
<output>
<ID>OUT_1</ID>272 </output>
<output>
<ID>OUT_2</ID>273 </output>
<output>
<ID>OUT_3</ID>274 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>214</ID>
<type>DD_KEYPAD_HEX</type>
<position>60,-38</position>
<output>
<ID>OUT_0</ID>275 </output>
<output>
<ID>OUT_1</ID>276 </output>
<output>
<ID>OUT_2</ID>277 </output>
<output>
<ID>OUT_3</ID>278 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>215</ID>
<type>BB_CLOCK</type>
<position>48.5,-75.5</position>
<output>
<ID>CLK</ID>330 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>77.5,-25</position>
<output>
<ID>OUT_0</ID>294 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>65,-27</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>65,-24.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_TOGGLE</type>
<position>90.5,-27.5</position>
<output>
<ID>OUT_0</ID>293 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>78.5,-72.5</position>
<output>
<ID>OUT_0</ID>310 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>73,-69.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_TOGGLE</type>
<position>129.5,-54</position>
<output>
<ID>OUT_0</ID>295 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>74.5,-36</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>91,-36</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>111.5,-35</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>133.5,-51</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_TOGGLE</type>
<position>146.5,-53.5</position>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>228</ID>
<type>BE_ROM_8x8</type>
<position>164.5,-61</position>
<input>
<ID>ADDRESS_0</ID>307 </input>
<input>
<ID>ADDRESS_1</ID>308 </input>
<input>
<ID>ENABLE_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_TOGGLE</type>
<position>121.5,-41</position>
<output>
<ID>OUT_0</ID>311 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_TOGGLE</type>
<position>121.5,-44</position>
<output>
<ID>OUT_0</ID>312 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>128,-40.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>128.5,-43.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>125.5,-61</position>
<input>
<ID>ENABLE_0</ID>312 </input>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>313 </input>
<input>
<ID>IN_2</ID>314 </input>
<input>
<ID>IN_3</ID>315 </input>
<input>
<ID>IN_4</ID>316 </input>
<input>
<ID>IN_5</ID>317 </input>
<input>
<ID>IN_6</ID>318 </input>
<input>
<ID>IN_7</ID>319 </input>
<output>
<ID>OUT_0</ID>321 </output>
<output>
<ID>OUT_1</ID>322 </output>
<output>
<ID>OUT_2</ID>323 </output>
<output>
<ID>OUT_3</ID>324 </output>
<output>
<ID>OUT_4</ID>325 </output>
<output>
<ID>OUT_5</ID>320 </output>
<output>
<ID>OUT_6</ID>327 </output>
<output>
<ID>OUT_7</ID>326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>234</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>104.5,-61</position>
<input>
<ID>ENABLE_0</ID>311 </input>
<output>
<ID>OUT_0</ID>328 </output>
<output>
<ID>OUT_1</ID>313 </output>
<output>
<ID>OUT_2</ID>314 </output>
<output>
<ID>OUT_3</ID>315 </output>
<output>
<ID>OUT_4</ID>316 </output>
<output>
<ID>OUT_5</ID>317 </output>
<output>
<ID>OUT_6</ID>318 </output>
<output>
<ID>OUT_7</ID>319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>151,-53</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>173.5,-61.5</position>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>175,-58.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AA_AND2</type>
<position>74.5,-57</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>332 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>60,-74.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_TOGGLE</type>
<position>54.5,-71.5</position>
<output>
<ID>OUT_0</ID>331 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_TOGGLE</type>
<position>45.5,-58</position>
<output>
<ID>OUT_0</ID>333 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>242</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>98.5,-116.5</position>
<input>
<ID>ENABLE_0</ID>354 </input>
<input>
<ID>IN_0</ID>335 </input>
<input>
<ID>IN_1</ID>336 </input>
<input>
<ID>IN_10</ID>345 </input>
<input>
<ID>IN_11</ID>346 </input>
<input>
<ID>IN_12</ID>347 </input>
<input>
<ID>IN_13</ID>348 </input>
<input>
<ID>IN_14</ID>349 </input>
<input>
<ID>IN_15</ID>350 </input>
<input>
<ID>IN_2</ID>337 </input>
<input>
<ID>IN_3</ID>338 </input>
<input>
<ID>IN_4</ID>339 </input>
<input>
<ID>IN_5</ID>340 </input>
<input>
<ID>IN_6</ID>341 </input>
<input>
<ID>IN_7</ID>342 </input>
<input>
<ID>IN_8</ID>343 </input>
<input>
<ID>IN_9</ID>344 </input>
<output>
<ID>OUT_0</ID>372 </output>
<output>
<ID>OUT_1</ID>373 </output>
<output>
<ID>OUT_10</ID>382 </output>
<output>
<ID>OUT_11</ID>383 </output>
<output>
<ID>OUT_12</ID>384 </output>
<output>
<ID>OUT_13</ID>385 </output>
<output>
<ID>OUT_14</ID>386 </output>
<output>
<ID>OUT_15</ID>387 </output>
<output>
<ID>OUT_2</ID>374 </output>
<output>
<ID>OUT_3</ID>375 </output>
<output>
<ID>OUT_4</ID>376 </output>
<output>
<ID>OUT_5</ID>377 </output>
<output>
<ID>OUT_6</ID>378 </output>
<output>
<ID>OUT_7</ID>379 </output>
<output>
<ID>OUT_8</ID>380 </output>
<output>
<ID>OUT_9</ID>381 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>243</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>98.5,-139.5</position>
<input>
<ID>ENABLE_0</ID>353 </input>
<input>
<ID>IN_0</ID>335 </input>
<input>
<ID>IN_1</ID>336 </input>
<input>
<ID>IN_10</ID>345 </input>
<input>
<ID>IN_11</ID>346 </input>
<input>
<ID>IN_12</ID>347 </input>
<input>
<ID>IN_13</ID>348 </input>
<input>
<ID>IN_14</ID>349 </input>
<input>
<ID>IN_15</ID>350 </input>
<input>
<ID>IN_2</ID>337 </input>
<input>
<ID>IN_3</ID>338 </input>
<input>
<ID>IN_4</ID>339 </input>
<input>
<ID>IN_5</ID>340 </input>
<input>
<ID>IN_6</ID>341 </input>
<input>
<ID>IN_7</ID>342 </input>
<input>
<ID>IN_8</ID>343 </input>
<input>
<ID>IN_9</ID>344 </input>
<output>
<ID>OUT_0</ID>356 </output>
<output>
<ID>OUT_1</ID>364 </output>
<output>
<ID>OUT_10</ID>361 </output>
<output>
<ID>OUT_11</ID>369 </output>
<output>
<ID>OUT_12</ID>362 </output>
<output>
<ID>OUT_13</ID>370 </output>
<output>
<ID>OUT_14</ID>363 </output>
<output>
<ID>OUT_15</ID>371 </output>
<output>
<ID>OUT_2</ID>357 </output>
<output>
<ID>OUT_3</ID>365 </output>
<output>
<ID>OUT_4</ID>358 </output>
<output>
<ID>OUT_5</ID>366 </output>
<output>
<ID>OUT_6</ID>359 </output>
<output>
<ID>OUT_7</ID>367 </output>
<output>
<ID>OUT_8</ID>360 </output>
<output>
<ID>OUT_9</ID>368 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>76,-103.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>DD_KEYPAD_HEX</type>
<position>58.5,-110</position>
<output>
<ID>OUT_0</ID>344 </output>
<output>
<ID>OUT_1</ID>346 </output>
<output>
<ID>OUT_2</ID>348 </output>
<output>
<ID>OUT_3</ID>350 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>246</ID>
<type>DD_KEYPAD_HEX</type>
<position>58.5,-134</position>
<output>
<ID>OUT_0</ID>343 </output>
<output>
<ID>OUT_1</ID>345 </output>
<output>
<ID>OUT_2</ID>347 </output>
<output>
<ID>OUT_3</ID>349 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>247</ID>
<type>DD_KEYPAD_HEX</type>
<position>58.5,-122</position>
<output>
<ID>OUT_0</ID>336 </output>
<output>
<ID>OUT_1</ID>338 </output>
<output>
<ID>OUT_2</ID>340 </output>
<output>
<ID>OUT_3</ID>342 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>248</ID>
<type>DD_KEYPAD_HEX</type>
<position>58.5,-146</position>
<output>
<ID>OUT_0</ID>335 </output>
<output>
<ID>OUT_1</ID>337 </output>
<output>
<ID>OUT_2</ID>339 </output>
<output>
<ID>OUT_3</ID>341 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_LABEL</type>
<position>49,-135</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>48.5,-109</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>48.5,-121.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>48.5,-146.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>BA_DECODER_2x4</type>
<position>90,-100</position>
<input>
<ID>ENABLE</ID>351 </input>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>353 </output>
<output>
<ID>OUT_1</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>85,-98.5</position>
<output>
<ID>OUT_0</ID>351 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>80.5,-101.5</position>
<output>
<ID>OUT_0</ID>352 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>85.5,-95.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>74,-101</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AE_FULLADDER_4BIT</type>
<position>116,-135.5</position>
<input>
<ID>IN_0</ID>364 </input>
<input>
<ID>IN_1</ID>365 </input>
<input>
<ID>IN_2</ID>366 </input>
<input>
<ID>IN_3</ID>367 </input>
<input>
<ID>IN_B_0</ID>356 </input>
<input>
<ID>IN_B_1</ID>357 </input>
<input>
<ID>IN_B_2</ID>358 </input>
<input>
<ID>IN_B_3</ID>359 </input>
<output>
<ID>OUT_0</ID>388 </output>
<output>
<ID>OUT_1</ID>389 </output>
<output>
<ID>OUT_2</ID>390 </output>
<output>
<ID>OUT_3</ID>391 </output>
<output>
<ID>carry_out</ID>355 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_FULLADDER_4BIT</type>
<position>116,-151.5</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>369 </input>
<input>
<ID>IN_2</ID>370 </input>
<input>
<ID>IN_3</ID>371 </input>
<input>
<ID>IN_B_0</ID>360 </input>
<input>
<ID>IN_B_1</ID>361 </input>
<input>
<ID>IN_B_2</ID>362 </input>
<input>
<ID>IN_B_3</ID>363 </input>
<output>
<ID>OUT_0</ID>392 </output>
<output>
<ID>OUT_1</ID>393 </output>
<output>
<ID>OUT_2</ID>394 </output>
<output>
<ID>OUT_3</ID>395 </output>
<input>
<ID>carry_in</ID>355 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>123.5,-128</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>124,-156.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>109.5,-129</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>110,-135.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>109.5,-145</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>110.5,-152</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_AND2</type>
<position>111.5,-125</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_AND2</type>
<position>116.5,-121.5</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>374 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>111.5,-118</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_AND2</type>
<position>116.5,-114.5</position>
<input>
<ID>IN_0</ID>379 </input>
<input>
<ID>IN_1</ID>378 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_AND2</type>
<position>111.5,-111</position>
<input>
<ID>IN_0</ID>381 </input>
<input>
<ID>IN_1</ID>380 </input>
<output>
<ID>OUT</ID>400 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>116.5,-107.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>382 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_AND2</type>
<position>111.5,-104</position>
<input>
<ID>IN_0</ID>385 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_AND2</type>
<position>116.5,-100.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>386 </input>
<output>
<ID>OUT</ID>403 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-112</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>403 </input>
<output>
<ID>OUT</ID>411 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-117</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>402 </input>
<output>
<ID>OUT</ID>410 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-122</position>
<input>
<ID>IN_0</ID>393 </input>
<input>
<ID>IN_1</ID>401 </input>
<output>
<ID>OUT</ID>409 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-127</position>
<input>
<ID>IN_0</ID>392 </input>
<input>
<ID>IN_1</ID>400 </input>
<output>
<ID>OUT</ID>408 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-132</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>399 </input>
<output>
<ID>OUT</ID>407 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-137</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>406 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-142</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>405 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_MUX_2x1</type>
<position>141.5,-147</position>
<input>
<ID>IN_0</ID>388 </input>
<input>
<ID>IN_1</ID>396 </input>
<output>
<ID>OUT</ID>404 </output>
<input>
<ID>SEL_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>164,-129</position>
<input>
<ID>IN_0</ID>404 </input>
<input>
<ID>IN_1</ID>405 </input>
<input>
<ID>IN_2</ID>406 </input>
<input>
<ID>IN_3</ID>407 </input>
<input>
<ID>IN_4</ID>408 </input>
<input>
<ID>IN_5</ID>409 </input>
<input>
<ID>IN_6</ID>410 </input>
<input>
<ID>IN_7</ID>411 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_LABEL</type>
<position>141.5,-150.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>142.5,-108</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>285</ID>
<type>GA_LED</type>
<position>155.5,-139</position>
<input>
<ID>N_in2</ID>411 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>286</ID>
<type>GA_LED</type>
<position>158,-139</position>
<input>
<ID>N_in2</ID>410 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>287</ID>
<type>GA_LED</type>
<position>160.5,-139</position>
<input>
<ID>N_in2</ID>409 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>288</ID>
<type>GA_LED</type>
<position>163,-139</position>
<input>
<ID>N_in2</ID>408 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>289</ID>
<type>GA_LED</type>
<position>165.5,-139</position>
<input>
<ID>N_in2</ID>407 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>290</ID>
<type>GA_LED</type>
<position>168,-139</position>
<input>
<ID>N_in2</ID>406 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>291</ID>
<type>GA_LED</type>
<position>170.5,-139</position>
<input>
<ID>N_in2</ID>405 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>292</ID>
<type>GA_LED</type>
<position>173,-139</position>
<input>
<ID>N_in2</ID>404 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>173,-141</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>170.5,-141</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_LABEL</type>
<position>168,-141</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_LABEL</type>
<position>165.5,-141</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>AA_LABEL</type>
<position>163,-141</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>298</ID>
<type>AA_LABEL</type>
<position>160.5,-141</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>AA_LABEL</type>
<position>158,-141</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>AA_LABEL</type>
<position>155.5,-141</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>AA_LABEL</type>
<position>291.5,-92.5</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AA_LABEL</type>
<position>291.5,-103.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>303</ID>
<type>AE_REGISTER8</type>
<position>234.5,-103.5</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>469 </input>
<input>
<ID>IN_4</ID>468 </input>
<input>
<ID>IN_5</ID>467 </input>
<input>
<ID>IN_6</ID>466 </input>
<input>
<ID>IN_7</ID>465 </input>
<output>
<ID>OUT_0</ID>435 </output>
<output>
<ID>OUT_1</ID>434 </output>
<output>
<ID>OUT_2</ID>433 </output>
<output>
<ID>OUT_3</ID>432 </output>
<output>
<ID>OUT_4</ID>431 </output>
<output>
<ID>OUT_5</ID>430 </output>
<output>
<ID>OUT_6</ID>429 </output>
<output>
<ID>OUT_7</ID>428 </output>
<input>
<ID>clock</ID>452 </input>
<input>
<ID>load</ID>475 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_REGISTER8</type>
<position>234.5,-116.5</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>469 </input>
<input>
<ID>IN_4</ID>468 </input>
<input>
<ID>IN_5</ID>467 </input>
<input>
<ID>IN_6</ID>466 </input>
<input>
<ID>IN_7</ID>465 </input>
<output>
<ID>OUT_0</ID>451 </output>
<output>
<ID>OUT_1</ID>442 </output>
<output>
<ID>OUT_2</ID>441 </output>
<output>
<ID>OUT_3</ID>440 </output>
<output>
<ID>OUT_4</ID>439 </output>
<output>
<ID>OUT_5</ID>438 </output>
<output>
<ID>OUT_6</ID>437 </output>
<output>
<ID>OUT_7</ID>436 </output>
<input>
<ID>clock</ID>452 </input>
<input>
<ID>load</ID>476 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>305</ID>
<type>AE_MUX_4x1</type>
<position>260,-66</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>428 </input>
<input>
<ID>IN_2</ID>420 </input>
<input>
<ID>IN_3</ID>412 </input>
<output>
<ID>OUT</ID>443 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_MUX_4x1</type>
<position>260,-77</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>429 </input>
<input>
<ID>IN_2</ID>421 </input>
<input>
<ID>IN_3</ID>413 </input>
<output>
<ID>OUT</ID>444 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_MUX_4x1</type>
<position>260,-88</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>430 </input>
<input>
<ID>IN_2</ID>422 </input>
<input>
<ID>IN_3</ID>414 </input>
<output>
<ID>OUT</ID>445 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_MUX_4x1</type>
<position>260,-97.5</position>
<input>
<ID>IN_0</ID>439 </input>
<input>
<ID>IN_1</ID>431 </input>
<input>
<ID>IN_2</ID>423 </input>
<input>
<ID>IN_3</ID>415 </input>
<output>
<ID>OUT</ID>446 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_MUX_4x1</type>
<position>260,-108.5</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>424 </input>
<input>
<ID>IN_3</ID>416 </input>
<output>
<ID>OUT</ID>447 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>310</ID>
<type>AE_MUX_4x1</type>
<position>260,-119.5</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>433 </input>
<input>
<ID>IN_2</ID>425 </input>
<input>
<ID>IN_3</ID>417 </input>
<output>
<ID>OUT</ID>448 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>209.5,-17.5</position>
<gparam>LABEL_TEXT Not most recent update</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AE_MUX_4x1</type>
<position>260,-130</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>434 </input>
<input>
<ID>IN_2</ID>426 </input>
<input>
<ID>IN_3</ID>418 </input>
<output>
<ID>OUT</ID>449 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_MUX_4x1</type>
<position>260,-141</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>435 </input>
<input>
<ID>IN_2</ID>427 </input>
<input>
<ID>IN_3</ID>419 </input>
<output>
<ID>OUT</ID>450 </output>
<input>
<ID>SEL_0</ID>453 </input>
<input>
<ID>SEL_1</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>313</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>292,-98.5</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>449 </input>
<input>
<ID>IN_2</ID>448 </input>
<input>
<ID>IN_3</ID>447 </input>
<input>
<ID>IN_4</ID>446 </input>
<input>
<ID>IN_5</ID>445 </input>
<input>
<ID>IN_6</ID>444 </input>
<input>
<ID>IN_7</ID>443 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>197,-31.5</position>
<gparam>LABEL_TEXT Check page 5</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>DD_KEYPAD_HEX</type>
<position>201.5,-81</position>
<output>
<ID>OUT_0</ID>453 </output>
<output>
<ID>OUT_1</ID>454 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>315</ID>
<type>BB_CLOCK</type>
<position>223,-125</position>
<output>
<ID>CLK</ID>452 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_LABEL</type>
<position>235.5,-70</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>AA_LABEL</type>
<position>235.5,-83</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>235.5,-96.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>AA_LABEL</type>
<position>235.5,-109.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AA_LABEL</type>
<position>200,-74</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>321</ID>
<type>DD_KEYPAD_HEX</type>
<position>201.5,-95</position>
<output>
<ID>OUT_0</ID>463 </output>
<output>
<ID>OUT_1</ID>464 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-66</position>
<input>
<ID>IN_0</ID>412 </input>
<input>
<ID>IN_1</ID>428 </input>
<input>
<ID>IN_2</ID>420 </input>
<input>
<ID>IN_3</ID>412 </input>
<output>
<ID>OUT</ID>455 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-77</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>429 </input>
<input>
<ID>IN_2</ID>421 </input>
<input>
<ID>IN_3</ID>413 </input>
<output>
<ID>OUT</ID>456 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-88</position>
<input>
<ID>IN_0</ID>438 </input>
<input>
<ID>IN_1</ID>430 </input>
<input>
<ID>IN_2</ID>422 </input>
<input>
<ID>IN_3</ID>414 </input>
<output>
<ID>OUT</ID>457 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>325</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-97.5</position>
<input>
<ID>IN_0</ID>439 </input>
<input>
<ID>IN_1</ID>431 </input>
<input>
<ID>IN_2</ID>423 </input>
<input>
<ID>IN_3</ID>415 </input>
<output>
<ID>OUT</ID>458 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-108.5</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>432 </input>
<input>
<ID>IN_2</ID>424 </input>
<input>
<ID>IN_3</ID>416 </input>
<output>
<ID>OUT</ID>459 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>327</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-119.5</position>
<input>
<ID>IN_0</ID>441 </input>
<input>
<ID>IN_1</ID>433 </input>
<input>
<ID>IN_2</ID>425 </input>
<input>
<ID>IN_3</ID>417 </input>
<output>
<ID>OUT</ID>460 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-130</position>
<input>
<ID>IN_0</ID>442 </input>
<input>
<ID>IN_1</ID>434 </input>
<input>
<ID>IN_2</ID>426 </input>
<input>
<ID>IN_3</ID>418 </input>
<output>
<ID>OUT</ID>461 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>329</ID>
<type>AE_MUX_4x1</type>
<position>272.5,-141</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>435 </input>
<input>
<ID>IN_2</ID>427 </input>
<input>
<ID>IN_3</ID>419 </input>
<output>
<ID>OUT</ID>462 </output>
<input>
<ID>SEL_0</ID>463 </input>
<input>
<ID>SEL_1</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>330</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>292,-109.5</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>461 </input>
<input>
<ID>IN_2</ID>460 </input>
<input>
<ID>IN_3</ID>459 </input>
<input>
<ID>IN_4</ID>458 </input>
<input>
<ID>IN_5</ID>457 </input>
<input>
<ID>IN_6</ID>456 </input>
<input>
<ID>IN_7</ID>455 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_LABEL</type>
<position>200,-88</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>DD_KEYPAD_HEX</type>
<position>217.5,-94.5</position>
<output>
<ID>OUT_0</ID>468 </output>
<output>
<ID>OUT_1</ID>467 </output>
<output>
<ID>OUT_2</ID>466 </output>
<output>
<ID>OUT_3</ID>465 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>333</ID>
<type>DD_KEYPAD_HEX</type>
<position>217.5,-106.5</position>
<output>
<ID>OUT_0</ID>472 </output>
<output>
<ID>OUT_1</ID>471 </output>
<output>
<ID>OUT_2</ID>470 </output>
<output>
<ID>OUT_3</ID>469 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_LABEL</type>
<position>217.5,-87.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>335</ID>
<type>BA_DECODER_2x4</type>
<position>219.5,-61.5</position>
<input>
<ID>ENABLE</ID>477 </input>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT_0</ID>473 </output>
<output>
<ID>OUT_1</ID>474 </output>
<output>
<ID>OUT_2</ID>475 </output>
<output>
<ID>OUT_3</ID>476 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_TOGGLE</type>
<position>213.5,-61</position>
<output>
<ID>OUT_0</ID>477 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_LABEL</type>
<position>211,-59.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>DD_KEYPAD_HEX</type>
<position>214.5,-74</position>
<output>
<ID>OUT_0</ID>478 </output>
<output>
<ID>OUT_1</ID>479 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>215,-67</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>AE_REGISTER8</type>
<position>234.5,-77</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>469 </input>
<input>
<ID>IN_4</ID>468 </input>
<input>
<ID>IN_5</ID>467 </input>
<input>
<ID>IN_6</ID>466 </input>
<input>
<ID>IN_7</ID>465 </input>
<output>
<ID>OUT_0</ID>419 </output>
<output>
<ID>OUT_1</ID>418 </output>
<output>
<ID>OUT_2</ID>417 </output>
<output>
<ID>OUT_3</ID>416 </output>
<output>
<ID>OUT_4</ID>415 </output>
<output>
<ID>OUT_5</ID>414 </output>
<output>
<ID>OUT_6</ID>413 </output>
<output>
<ID>OUT_7</ID>412 </output>
<input>
<ID>clock</ID>452 </input>
<input>
<ID>load</ID>473 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>341</ID>
<type>AE_REGISTER8</type>
<position>234.5,-90</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>470 </input>
<input>
<ID>IN_3</ID>469 </input>
<input>
<ID>IN_4</ID>468 </input>
<input>
<ID>IN_5</ID>467 </input>
<input>
<ID>IN_6</ID>466 </input>
<input>
<ID>IN_7</ID>465 </input>
<output>
<ID>OUT_0</ID>427 </output>
<output>
<ID>OUT_1</ID>426 </output>
<output>
<ID>OUT_2</ID>425 </output>
<output>
<ID>OUT_3</ID>424 </output>
<output>
<ID>OUT_4</ID>423 </output>
<output>
<ID>OUT_5</ID>422 </output>
<output>
<ID>OUT_6</ID>421 </output>
<output>
<ID>OUT_7</ID>420 </output>
<input>
<ID>clock</ID>452 </input>
<input>
<ID>load</ID>474 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>245,-52.5</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-143,129.5,-135</points>
<intersection>-143 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-143,139.5,-143</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-135,129.5,-135</points>
<connection>
<GID>258</GID>
<name>OUT_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-138,129.5,-136</points>
<intersection>-138 1</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-138,139.5,-138</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-136,129.5,-136</points>
<connection>
<GID>258</GID>
<name>OUT_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-137,129.5,-133</points>
<intersection>-137 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-133,139.5,-133</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-137,129.5,-137</points>
<connection>
<GID>258</GID>
<name>OUT_3</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-150,129.5,-128</points>
<intersection>-150 2</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-128,139.5,-128</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-150,129.5,-150</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-151,129.5,-123</points>
<intersection>-151 2</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-123,139.5,-123</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-151,129.5,-151</points>
<connection>
<GID>259</GID>
<name>OUT_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-152,129.5,-118</points>
<intersection>-152 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-118,139.5,-118</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-152,129.5,-152</points>
<connection>
<GID>259</GID>
<name>OUT_2</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-153,129.5,-113</points>
<intersection>-153 2</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-113,139.5,-113</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-153,129.5,-153</points>
<connection>
<GID>259</GID>
<name>OUT_3</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-146,127,-125</points>
<intersection>-146 1</intersection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-146,139.5,-146</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-125,127,-125</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-141,129.5,-121.5</points>
<intersection>-141 2</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-121.5,129.5,-121.5</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-141,139.5,-141</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-136,127,-118</points>
<intersection>-136 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-118,127,-118</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-136,139.5,-136</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-131,129.5,-114.5</points>
<intersection>-131 2</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-114.5,129.5,-114.5</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-131,139.5,-131</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-126,127,-111</points>
<intersection>-126 2</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-111,127,-111</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-126,139.5,-126</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-121,129.5,-107.5</points>
<intersection>-121 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-107.5,129.5,-107.5</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-121,139.5,-121</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-116,127,-104</points>
<intersection>-116 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-104,127,-104</points>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-116,139.5,-116</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-111,129.5,-100.5</points>
<intersection>-111 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-100.5,129.5,-100.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-111,139.5,-111</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-147,151,-132</points>
<intersection>-147 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-132,159,-132</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection>
<intersection>152 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-147,151,-147</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>152,-137.5,152,-132</points>
<intersection>-137.5 8</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>152,-137.5,173,-137.5</points>
<intersection>152 7</intersection>
<intersection>173 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>173,-138,173,-137.5</points>
<connection>
<GID>292</GID>
<name>N_in2</name></connection>
<intersection>-137.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-142,151,-131</points>
<intersection>-142 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-131,159,-131</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection>
<intersection>152.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-142,151,-142</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>152.5,-137,152.5,-131</points>
<intersection>-137 8</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>152.5,-137,170.5,-137</points>
<intersection>152.5 7</intersection>
<intersection>170.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>170.5,-138,170.5,-137</points>
<connection>
<GID>291</GID>
<name>N_in2</name></connection>
<intersection>-137 8</intersection></vsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-137,151,-130</points>
<intersection>-137 2</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-130,159,-130</points>
<connection>
<GID>282</GID>
<name>IN_2</name></connection>
<intersection>151 0</intersection>
<intersection>153 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-137,151,-137</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>153,-136.5,153,-130</points>
<intersection>-136.5 8</intersection>
<intersection>-130 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>153,-136.5,168,-136.5</points>
<intersection>153 7</intersection>
<intersection>168 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>168,-138,168,-136.5</points>
<connection>
<GID>290</GID>
<name>N_in2</name></connection>
<intersection>-136.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-132,151,-129</points>
<intersection>-132 2</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-129,159,-129</points>
<connection>
<GID>282</GID>
<name>IN_3</name></connection>
<intersection>151 0</intersection>
<intersection>153.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-132,151,-132</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>153.5,-136,153.5,-129</points>
<intersection>-136 9</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>153.5,-136,165.5,-136</points>
<intersection>153.5 8</intersection>
<intersection>165.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>165.5,-138,165.5,-136</points>
<connection>
<GID>289</GID>
<name>N_in2</name></connection>
<intersection>-136 9</intersection></vsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-128,151,-127</points>
<intersection>-128 1</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-128,159,-128</points>
<connection>
<GID>282</GID>
<name>IN_4</name></connection>
<intersection>151 0</intersection>
<intersection>154 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-127,151,-127</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>154,-135.5,154,-128</points>
<intersection>-135.5 9</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>154,-135.5,163,-135.5</points>
<intersection>154 8</intersection>
<intersection>163 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>163,-138,163,-135.5</points>
<connection>
<GID>288</GID>
<name>N_in2</name></connection>
<intersection>-135.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-127,151,-122</points>
<intersection>-127 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-127,159,-127</points>
<connection>
<GID>282</GID>
<name>IN_5</name></connection>
<intersection>151 0</intersection>
<intersection>154.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-122,151,-122</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>154.5,-135,154.5,-127</points>
<intersection>-135 8</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>154.5,-135,160.5,-135</points>
<intersection>154.5 7</intersection>
<intersection>160.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>160.5,-138,160.5,-135</points>
<connection>
<GID>287</GID>
<name>N_in2</name></connection>
<intersection>-135 8</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-126,151,-117</points>
<intersection>-126 1</intersection>
<intersection>-117 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-126,159,-126</points>
<connection>
<GID>282</GID>
<name>IN_6</name></connection>
<intersection>151 0</intersection>
<intersection>155 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-117,151,-117</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>155,-134.5,155,-126</points>
<intersection>-134.5 8</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>155,-134.5,158,-134.5</points>
<intersection>155 7</intersection>
<intersection>158 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>158,-138,158,-134.5</points>
<connection>
<GID>286</GID>
<name>N_in2</name></connection>
<intersection>-134.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-125,151,-112</points>
<intersection>-125 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,-112,151,-112</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-125,159,-125</points>
<connection>
<GID>282</GID>
<name>IN_7</name></connection>
<intersection>151 0</intersection>
<intersection>155.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>155.5,-138,155.5,-125</points>
<connection>
<GID>285</GID>
<name>N_in2</name></connection>
<intersection>-125 2</intersection></vsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-73,256.5,-73</points>
<connection>
<GID>340</GID>
<name>OUT_7</name></connection>
<intersection>256.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>256.5,-73,256.5,-63</points>
<intersection>-73 1</intersection>
<intersection>-63 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>256.5,-63,269.5,-63</points>
<connection>
<GID>305</GID>
<name>IN_3</name></connection>
<connection>
<GID>322</GID>
<name>IN_3</name></connection>
<intersection>256.5 4</intersection>
<intersection>268 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>268,-69,268,-63</points>
<intersection>-69 8</intersection>
<intersection>-63 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>268,-69,269.5,-69</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>268 6</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-74,269.5,-74</points>
<connection>
<GID>340</GID>
<name>OUT_6</name></connection>
<connection>
<GID>323</GID>
<name>IN_3</name></connection>
<connection>
<GID>306</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-85,255.5,-75</points>
<intersection>-85 1</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-85,269.5,-85</points>
<connection>
<GID>307</GID>
<name>IN_3</name></connection>
<connection>
<GID>324</GID>
<name>IN_3</name></connection>
<intersection>255.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-75,255.5,-75</points>
<connection>
<GID>340</GID>
<name>OUT_5</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-94.5,255,-76</points>
<intersection>-94.5 1</intersection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,-94.5,269.5,-94.5</points>
<connection>
<GID>308</GID>
<name>IN_3</name></connection>
<connection>
<GID>325</GID>
<name>IN_3</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-76,255,-76</points>
<connection>
<GID>340</GID>
<name>OUT_4</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-105.5,254.5,-77</points>
<intersection>-105.5 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254.5,-105.5,269.5,-105.5</points>
<connection>
<GID>309</GID>
<name>IN_3</name></connection>
<connection>
<GID>326</GID>
<name>IN_3</name></connection>
<intersection>254.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-77,254.5,-77</points>
<connection>
<GID>340</GID>
<name>OUT_3</name></connection>
<intersection>254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254,-116.5,254,-78</points>
<intersection>-116.5 1</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254,-116.5,269.5,-116.5</points>
<connection>
<GID>310</GID>
<name>IN_3</name></connection>
<connection>
<GID>327</GID>
<name>IN_3</name></connection>
<intersection>254 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-78,254,-78</points>
<connection>
<GID>340</GID>
<name>OUT_2</name></connection>
<intersection>254 0</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253.5,-127,253.5,-79</points>
<intersection>-127 1</intersection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253.5,-127,269.5,-127</points>
<connection>
<GID>311</GID>
<name>IN_3</name></connection>
<connection>
<GID>328</GID>
<name>IN_3</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-79,253.5,-79</points>
<connection>
<GID>340</GID>
<name>OUT_1</name></connection>
<intersection>253.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253,-138,253,-80</points>
<intersection>-138 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,-80,253,-80</points>
<connection>
<GID>340</GID>
<name>OUT_0</name></connection>
<intersection>253 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>253,-138,269.5,-138</points>
<connection>
<GID>312</GID>
<name>IN_3</name></connection>
<connection>
<GID>329</GID>
<name>IN_3</name></connection>
<intersection>253 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252,-86,252,-65</points>
<intersection>-86 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252,-65,269.5,-65</points>
<connection>
<GID>305</GID>
<name>IN_2</name></connection>
<connection>
<GID>322</GID>
<name>IN_2</name></connection>
<intersection>252 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-86,252,-86</points>
<connection>
<GID>341</GID>
<name>OUT_7</name></connection>
<intersection>252 0</intersection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,-87,251.5,-76</points>
<intersection>-87 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251.5,-76,269.5,-76</points>
<connection>
<GID>306</GID>
<name>IN_2</name></connection>
<connection>
<GID>323</GID>
<name>IN_2</name></connection>
<intersection>251.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-87,251.5,-87</points>
<connection>
<GID>341</GID>
<name>OUT_6</name></connection>
<intersection>251.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-88,257,-88</points>
<connection>
<GID>341</GID>
<name>OUT_5</name></connection>
<intersection>257 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>257,-88,257,-87</points>
<connection>
<GID>307</GID>
<name>IN_2</name></connection>
<intersection>-88 1</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>257,-87,269.5,-87</points>
<connection>
<GID>324</GID>
<name>IN_2</name></connection>
<intersection>257 3</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-96.5,251,-89</points>
<intersection>-96.5 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,-96.5,269.5,-96.5</points>
<connection>
<GID>308</GID>
<name>IN_2</name></connection>
<connection>
<GID>325</GID>
<name>IN_2</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-89,251,-89</points>
<connection>
<GID>341</GID>
<name>OUT_4</name></connection>
<intersection>251 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,-107.5,250.5,-90</points>
<intersection>-107.5 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,-107.5,269.5,-107.5</points>
<connection>
<GID>309</GID>
<name>IN_2</name></connection>
<connection>
<GID>326</GID>
<name>IN_2</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-90,250.5,-90</points>
<connection>
<GID>341</GID>
<name>OUT_3</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-118.5,250,-91</points>
<intersection>-118.5 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,-118.5,269.5,-118.5</points>
<connection>
<GID>310</GID>
<name>IN_2</name></connection>
<connection>
<GID>327</GID>
<name>IN_2</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-91,250,-91</points>
<connection>
<GID>341</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-129,249.5,-92</points>
<intersection>-129 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,-92,249.5,-92</points>
<connection>
<GID>341</GID>
<name>OUT_1</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-129,269.5,-129</points>
<connection>
<GID>311</GID>
<name>IN_2</name></connection>
<connection>
<GID>328</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,-140,252.5,-93</points>
<intersection>-140 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252.5,-140,269.5,-140</points>
<connection>
<GID>312</GID>
<name>IN_2</name></connection>
<connection>
<GID>329</GID>
<name>IN_2</name></connection>
<intersection>252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-93,252.5,-93</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-99.5,248,-67</points>
<intersection>-99.5 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-67,269.5,-67</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-99.5,248,-99.5</points>
<connection>
<GID>303</GID>
<name>OUT_7</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,-100.5,247.5,-78</points>
<intersection>-100.5 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,-78,269.5,-78</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-100.5,247.5,-100.5</points>
<connection>
<GID>303</GID>
<name>OUT_6</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,-101.5,247,-89</points>
<intersection>-101.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,-89,269.5,-89</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-101.5,247,-101.5</points>
<connection>
<GID>303</GID>
<name>OUT_5</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-102.5,246.5,-98.5</points>
<intersection>-102.5 2</intersection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246.5,-98.5,269.5,-98.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-102.5,246.5,-102.5</points>
<connection>
<GID>303</GID>
<name>OUT_4</name></connection>
<intersection>246.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-109.5,246,-103.5</points>
<intersection>-109.5 1</intersection>
<intersection>-103.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246,-109.5,269.5,-109.5</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-103.5,246,-103.5</points>
<connection>
<GID>303</GID>
<name>OUT_3</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-120.5,245.5,-104.5</points>
<intersection>-120.5 1</intersection>
<intersection>-104.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-120.5,269.5,-120.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-104.5,245.5,-104.5</points>
<connection>
<GID>303</GID>
<name>OUT_2</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-131,245,-105.5</points>
<intersection>-131 1</intersection>
<intersection>-105.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-131,269.5,-131</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-105.5,245,-105.5</points>
<connection>
<GID>303</GID>
<name>OUT_1</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-142,244.5,-106.5</points>
<intersection>-142 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238.5,-106.5,244.5,-106.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244.5,-142,269.5,-142</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243.5,-112.5,243.5,-69</points>
<intersection>-112.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243.5,-69,257,-69</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>243.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-112.5,243.5,-112.5</points>
<connection>
<GID>304</GID>
<name>OUT_7</name></connection>
<intersection>243.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-113.5,243,-80</points>
<intersection>-113.5 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-80,269.5,-80</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-113.5,243,-113.5</points>
<connection>
<GID>304</GID>
<name>OUT_6</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-114.5,242.5,-91</points>
<intersection>-114.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>242.5,-91,269.5,-91</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>242.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-114.5,242.5,-114.5</points>
<connection>
<GID>304</GID>
<name>OUT_5</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>238.5,-100.5,269.5,-100.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>238.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>238.5,-115.5,238.5,-100.5</points>
<connection>
<GID>304</GID>
<name>OUT_4</name></connection>
<intersection>-100.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-116.5,241.5,-111.5</points>
<intersection>-116.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241.5,-111.5,269.5,-111.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>241.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-116.5,241.5,-116.5</points>
<connection>
<GID>304</GID>
<name>OUT_3</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-122.5,241,-117.5</points>
<intersection>-122.5 1</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-122.5,269.5,-122.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>241 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-117.5,241,-117.5</points>
<connection>
<GID>304</GID>
<name>OUT_2</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-133,240.5,-118.5</points>
<intersection>-133 1</intersection>
<intersection>-118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240.5,-133,269.5,-133</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>240.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-118.5,240.5,-118.5</points>
<connection>
<GID>304</GID>
<name>OUT_1</name></connection>
<intersection>240.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-94.5,281.5,-66</points>
<intersection>-94.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-66,281.5,-66</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-94.5,287,-94.5</points>
<connection>
<GID>313</GID>
<name>IN_7</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-95.5,281.5,-77</points>
<intersection>-95.5 2</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-77,281.5,-77</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-95.5,287,-95.5</points>
<connection>
<GID>313</GID>
<name>IN_6</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-96.5,281.5,-88</points>
<intersection>-96.5 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-88,281.5,-88</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-96.5,287,-96.5</points>
<connection>
<GID>313</GID>
<name>IN_5</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>263,-97.5,287,-97.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<connection>
<GID>313</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-108.5,281.5,-98.5</points>
<intersection>-108.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-108.5,281.5,-108.5</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-98.5,287,-98.5</points>
<connection>
<GID>313</GID>
<name>IN_3</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-119.5,281.5,-99.5</points>
<intersection>-119.5 1</intersection>
<intersection>-99.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-119.5,281.5,-119.5</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-99.5,287,-99.5</points>
<connection>
<GID>313</GID>
<name>IN_2</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-130,281.5,-100.5</points>
<intersection>-130 1</intersection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-130,281.5,-130</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-100.5,287,-100.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-141,281.5,-101.5</points>
<intersection>-141 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-101.5,287,-101.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>263,-141,281.5,-141</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-144,240,-119.5</points>
<intersection>-144 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-144,269.5,-144</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>238.5,-119.5,240,-119.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,-125,230,-82</points>
<intersection>-125 10</intersection>
<intersection>-121.5 8</intersection>
<intersection>-108.5 7</intersection>
<intersection>-95 6</intersection>
<intersection>-82 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>230,-82,233.5,-82</points>
<connection>
<GID>340</GID>
<name>clock</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>230,-95,233.5,-95</points>
<connection>
<GID>341</GID>
<name>clock</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>230,-108.5,233.5,-108.5</points>
<connection>
<GID>303</GID>
<name>clock</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>230,-121.5,233.5,-121.5</points>
<connection>
<GID>304</GID>
<name>clock</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>227,-125,230,-125</points>
<connection>
<GID>315</GID>
<name>CLK</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261,-136,261,-58</points>
<connection>
<GID>312</GID>
<name>SEL_0</name></connection>
<connection>
<GID>311</GID>
<name>SEL_0</name></connection>
<connection>
<GID>310</GID>
<name>SEL_0</name></connection>
<connection>
<GID>309</GID>
<name>SEL_0</name></connection>
<connection>
<GID>308</GID>
<name>SEL_0</name></connection>
<connection>
<GID>307</GID>
<name>SEL_0</name></connection>
<connection>
<GID>306</GID>
<name>SEL_0</name></connection>
<connection>
<GID>305</GID>
<name>SEL_0</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-58,261,-58</points>
<intersection>207.5 2</intersection>
<intersection>261 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>207.5,-84,207.5,-58</points>
<intersection>-84 3</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>206.5,-84,207.5,-84</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>207.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-136,260,-58.5</points>
<connection>
<GID>312</GID>
<name>SEL_1</name></connection>
<connection>
<GID>311</GID>
<name>SEL_1</name></connection>
<connection>
<GID>310</GID>
<name>SEL_1</name></connection>
<connection>
<GID>309</GID>
<name>SEL_1</name></connection>
<connection>
<GID>308</GID>
<name>SEL_1</name></connection>
<connection>
<GID>307</GID>
<name>SEL_1</name></connection>
<connection>
<GID>306</GID>
<name>SEL_1</name></connection>
<connection>
<GID>305</GID>
<name>SEL_1</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-58.5,260,-58.5</points>
<intersection>207 2</intersection>
<intersection>260 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>207,-82,207,-58.5</points>
<intersection>-82 3</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>206.5,-82,207,-82</points>
<connection>
<GID>314</GID>
<name>OUT_1</name></connection>
<intersection>207 2</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-105.5,276,-66</points>
<intersection>-105.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-66,276,-66</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-105.5,287,-105.5</points>
<connection>
<GID>330</GID>
<name>IN_7</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-106.5,276,-77</points>
<intersection>-106.5 2</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-77,276,-77</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-106.5,287,-106.5</points>
<connection>
<GID>330</GID>
<name>IN_6</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-107.5,276,-88</points>
<intersection>-107.5 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-88,276,-88</points>
<connection>
<GID>324</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-107.5,287,-107.5</points>
<connection>
<GID>330</GID>
<name>IN_5</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-108.5,276,-97.5</points>
<intersection>-108.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-97.5,276,-97.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-108.5,287,-108.5</points>
<connection>
<GID>330</GID>
<name>IN_4</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>276,-109.5,287,-109.5</points>
<connection>
<GID>330</GID>
<name>IN_3</name></connection>
<intersection>276 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>276,-109.5,276,-108.5</points>
<intersection>-109.5 1</intersection>
<intersection>-108.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>275.5,-108.5,276,-108.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>276 2</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-119.5,276,-110.5</points>
<intersection>-119.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-119.5,276,-119.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-110.5,287,-110.5</points>
<connection>
<GID>330</GID>
<name>IN_2</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-130,276,-111.5</points>
<intersection>-130 1</intersection>
<intersection>-111.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-130,276,-130</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-111.5,287,-111.5</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-141,276,-112.5</points>
<intersection>-141 2</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-112.5,287,-112.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>275.5,-141,276,-141</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-136,273.5,-59.5</points>
<connection>
<GID>329</GID>
<name>SEL_0</name></connection>
<connection>
<GID>328</GID>
<name>SEL_0</name></connection>
<connection>
<GID>327</GID>
<name>SEL_0</name></connection>
<connection>
<GID>326</GID>
<name>SEL_0</name></connection>
<connection>
<GID>325</GID>
<name>SEL_0</name></connection>
<connection>
<GID>324</GID>
<name>SEL_0</name></connection>
<connection>
<GID>323</GID>
<name>SEL_0</name></connection>
<connection>
<GID>322</GID>
<name>SEL_0</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-59.5,273.5,-59.5</points>
<intersection>208.5 2</intersection>
<intersection>273.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>208.5,-98,208.5,-59.5</points>
<intersection>-98 3</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>206.5,-98,208.5,-98</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>208.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-136,272.5,-59</points>
<connection>
<GID>329</GID>
<name>SEL_1</name></connection>
<connection>
<GID>328</GID>
<name>SEL_1</name></connection>
<connection>
<GID>327</GID>
<name>SEL_1</name></connection>
<connection>
<GID>326</GID>
<name>SEL_1</name></connection>
<connection>
<GID>325</GID>
<name>SEL_1</name></connection>
<connection>
<GID>324</GID>
<name>SEL_1</name></connection>
<connection>
<GID>323</GID>
<name>SEL_1</name></connection>
<connection>
<GID>322</GID>
<name>SEL_1</name></connection>
<intersection>-59 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>208,-59,272.5,-59</points>
<intersection>208 16</intersection>
<intersection>272.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>208,-96,208,-59</points>
<intersection>-96 18</intersection>
<intersection>-59 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>206.5,-96,208,-96</points>
<connection>
<GID>321</GID>
<name>OUT_1</name></connection>
<intersection>208 16</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-112.5,229,-73</points>
<intersection>-112.5 6</intersection>
<intersection>-99.5 3</intersection>
<intersection>-91.5 4</intersection>
<intersection>-86 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229,-73,230.5,-73</points>
<connection>
<GID>340</GID>
<name>IN_7</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>229,-86,230.5,-86</points>
<connection>
<GID>341</GID>
<name>IN_7</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>229,-99.5,230.5,-99.5</points>
<connection>
<GID>303</GID>
<name>IN_7</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>222.5,-91.5,229,-91.5</points>
<connection>
<GID>332</GID>
<name>OUT_3</name></connection>
<intersection>229 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>229,-112.5,230.5,-112.5</points>
<connection>
<GID>304</GID>
<name>IN_7</name></connection>
<intersection>229 0</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-113.5,228.5,-74</points>
<intersection>-113.5 6</intersection>
<intersection>-100.5 5</intersection>
<intersection>-93.5 2</intersection>
<intersection>-87 3</intersection>
<intersection>-74 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-93.5,228.5,-93.5</points>
<connection>
<GID>332</GID>
<name>OUT_2</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,-87,230.5,-87</points>
<connection>
<GID>341</GID>
<name>IN_6</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>228.5,-74,230.5,-74</points>
<connection>
<GID>340</GID>
<name>IN_6</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228.5,-100.5,230.5,-100.5</points>
<connection>
<GID>303</GID>
<name>IN_6</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228.5,-113.5,230.5,-113.5</points>
<connection>
<GID>304</GID>
<name>IN_6</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-114.5,228,-75</points>
<intersection>-114.5 6</intersection>
<intersection>-101.5 3</intersection>
<intersection>-95.5 2</intersection>
<intersection>-88 4</intersection>
<intersection>-75 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-95.5,228,-95.5</points>
<connection>
<GID>332</GID>
<name>OUT_1</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228,-101.5,230.5,-101.5</points>
<connection>
<GID>303</GID>
<name>IN_5</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>228,-88,230.5,-88</points>
<connection>
<GID>341</GID>
<name>IN_5</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>228,-75,230.5,-75</points>
<connection>
<GID>340</GID>
<name>IN_5</name></connection>
<intersection>228 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>228,-114.5,230.5,-114.5</points>
<connection>
<GID>304</GID>
<name>IN_5</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,-115.5,227.5,-76</points>
<intersection>-115.5 6</intersection>
<intersection>-102.5 3</intersection>
<intersection>-97.5 2</intersection>
<intersection>-89 4</intersection>
<intersection>-76 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-97.5,227.5,-97.5</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227.5,-102.5,230.5,-102.5</points>
<connection>
<GID>303</GID>
<name>IN_4</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>227.5,-89,230.5,-89</points>
<connection>
<GID>341</GID>
<name>IN_4</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227.5,-76,230.5,-76</points>
<connection>
<GID>340</GID>
<name>IN_4</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>227.5,-115.5,230.5,-115.5</points>
<connection>
<GID>304</GID>
<name>IN_4</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-116.5,227,-77</points>
<intersection>-116.5 5</intersection>
<intersection>-103.5 2</intersection>
<intersection>-90 3</intersection>
<intersection>-77 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-103.5,230.5,-103.5</points>
<connection>
<GID>303</GID>
<name>IN_3</name></connection>
<connection>
<GID>333</GID>
<name>OUT_3</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>227,-90,230.5,-90</points>
<connection>
<GID>341</GID>
<name>IN_3</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>227,-77,230.5,-77</points>
<connection>
<GID>340</GID>
<name>IN_3</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>227,-116.5,230.5,-116.5</points>
<connection>
<GID>304</GID>
<name>IN_3</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-117.5,226.5,-78</points>
<intersection>-117.5 5</intersection>
<intersection>-105.5 2</intersection>
<intersection>-104.5 4</intersection>
<intersection>-91 3</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,-78,230.5,-78</points>
<connection>
<GID>340</GID>
<name>IN_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-105.5,226.5,-105.5</points>
<connection>
<GID>333</GID>
<name>OUT_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>226.5,-91,230.5,-91</points>
<connection>
<GID>341</GID>
<name>IN_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226.5,-104.5,230.5,-104.5</points>
<connection>
<GID>303</GID>
<name>IN_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>226.5,-117.5,230.5,-117.5</points>
<connection>
<GID>304</GID>
<name>IN_2</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,-118.5,226,-79</points>
<intersection>-118.5 5</intersection>
<intersection>-107.5 2</intersection>
<intersection>-105.5 4</intersection>
<intersection>-92 3</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,-79,230.5,-79</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-107.5,226,-107.5</points>
<connection>
<GID>333</GID>
<name>OUT_1</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>226,-92,230.5,-92</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>226,-105.5,230.5,-105.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>226,-118.5,230.5,-118.5</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-119.5,225.5,-80</points>
<intersection>-119.5 5</intersection>
<intersection>-109.5 2</intersection>
<intersection>-106.5 4</intersection>
<intersection>-93 3</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-80,230.5,-80</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-109.5,225.5,-109.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>225.5,-93,230.5,-93</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>225.5,-106.5,230.5,-106.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-119.5,230.5,-119.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-71,232.5,-63</points>
<intersection>-71 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-63,232.5,-63</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232.5,-71,233.5,-71</points>
<connection>
<GID>340</GID>
<name>load</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-84,232.5,-62</points>
<intersection>-84 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-62,232.5,-62</points>
<connection>
<GID>335</GID>
<name>OUT_1</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232.5,-84,233.5,-84</points>
<connection>
<GID>341</GID>
<name>load</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-97.5,232.5,-61</points>
<intersection>-97.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-61,232.5,-61</points>
<connection>
<GID>335</GID>
<name>OUT_2</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232.5,-97.5,233.5,-97.5</points>
<connection>
<GID>303</GID>
<name>load</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-110.5,232.5,-60</points>
<intersection>-110.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-60,232.5,-60</points>
<connection>
<GID>335</GID>
<name>OUT_3</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>232.5,-110.5,233.5,-110.5</points>
<connection>
<GID>304</GID>
<name>load</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215.5,-61,216.5,-61</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>216.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>216.5,-61,216.5,-60</points>
<connection>
<GID>335</GID>
<name>ENABLE</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221,-77,221,-66</points>
<intersection>-77 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,-66,221,-66</points>
<intersection>216 3</intersection>
<intersection>221 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>219.5,-77,221,-77</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>221 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>216,-66,216,-63</points>
<intersection>-66 1</intersection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>216,-63,216.5,-63</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>216 3</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,-75,221.5,-65.5</points>
<intersection>-75 2</intersection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216.5,-65.5,221.5,-65.5</points>
<intersection>216.5 3</intersection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>219.5,-75,221.5,-75</points>
<connection>
<GID>338</GID>
<name>OUT_1</name></connection>
<intersection>221.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>216.5,-65.5,216.5,-62</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>-65.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-53,70,-47</points>
<intersection>-53 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-47,75.5,-47</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-53,70,-53</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-51,70,-46</points>
<intersection>-51 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-46,75.5,-46</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-51,70,-51</points>
<connection>
<GID>213</GID>
<name>OUT_1</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-49,70,-45</points>
<intersection>-49 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-45,75.5,-45</points>
<connection>
<GID>208</GID>
<name>IN_2</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-49,70,-49</points>
<connection>
<GID>213</GID>
<name>OUT_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-47,70,-44</points>
<intersection>-47 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-44,75.5,-44</points>
<connection>
<GID>208</GID>
<name>IN_3</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-47,70,-47</points>
<connection>
<GID>213</GID>
<name>OUT_3</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-43,70,-41</points>
<intersection>-43 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-43,75.5,-43</points>
<connection>
<GID>208</GID>
<name>IN_4</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-41,70,-41</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-42,70,-39</points>
<intersection>-42 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-42,75.5,-42</points>
<connection>
<GID>208</GID>
<name>IN_5</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-39,70,-39</points>
<connection>
<GID>214</GID>
<name>OUT_1</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-41,70,-37</points>
<intersection>-41 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-41,75.5,-41</points>
<connection>
<GID>208</GID>
<name>IN_6</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-37,70,-37</points>
<connection>
<GID>214</GID>
<name>OUT_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-40,75.5,-40</points>
<connection>
<GID>208</GID>
<name>IN_7</name></connection>
<intersection>65 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,-40,65,-35</points>
<connection>
<GID>214</GID>
<name>OUT_3</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-40,92.5,-40</points>
<connection>
<GID>209</GID>
<name>IN_7</name></connection>
<connection>
<GID>208</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-41,92.5,-41</points>
<connection>
<GID>209</GID>
<name>IN_6</name></connection>
<connection>
<GID>208</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-42,92.5,-42</points>
<connection>
<GID>209</GID>
<name>IN_5</name></connection>
<connection>
<GID>208</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-43,92.5,-43</points>
<connection>
<GID>209</GID>
<name>IN_4</name></connection>
<connection>
<GID>208</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-44,92.5,-44</points>
<connection>
<GID>209</GID>
<name>IN_3</name></connection>
<connection>
<GID>208</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-45,92.5,-45</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<connection>
<GID>208</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-46,92.5,-46</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<connection>
<GID>208</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,-47,92.5,-47</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-40,106.5,-40</points>
<connection>
<GID>211</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>209</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-41,106.5,-41</points>
<connection>
<GID>211</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>209</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-42,106.5,-42</points>
<connection>
<GID>211</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>209</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-43,106.5,-43</points>
<connection>
<GID>211</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>209</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-44,106.5,-44</points>
<connection>
<GID>211</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>209</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-45,106.5,-45</points>
<connection>
<GID>211</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>209</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-38,95.5,-27.5</points>
<connection>
<GID>209</GID>
<name>load</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-27.5,95.5,-27.5</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-38,79.5,-25</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<connection>
<GID>208</GID>
<name>count_enable</name></connection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-37,80.5,-37</points>
<intersection>79.5 0</intersection>
<intersection>80.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80.5,-38,80.5,-37</points>
<connection>
<GID>208</GID>
<name>count_up</name></connection>
<intersection>-37 2</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>131.5,-54,132.5,-54</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>132.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132.5,-55.5,132.5,-54</points>
<connection>
<GID>210</GID>
<name>load</name></connection>
<intersection>-54 2</intersection></vsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-46,106.5,-46</points>
<connection>
<GID>211</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>209</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-47,106.5,-47</points>
<connection>
<GID>211</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-57.5,145.5,-57.5</points>
<connection>
<GID>212</GID>
<name>IN_7</name></connection>
<connection>
<GID>210</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-58.5,145.5,-58.5</points>
<connection>
<GID>212</GID>
<name>IN_6</name></connection>
<connection>
<GID>210</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-59.5,145.5,-59.5</points>
<connection>
<GID>212</GID>
<name>IN_5</name></connection>
<connection>
<GID>210</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-60.5,145.5,-60.5</points>
<connection>
<GID>212</GID>
<name>IN_4</name></connection>
<connection>
<GID>210</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-61.5,145.5,-61.5</points>
<connection>
<GID>212</GID>
<name>IN_3</name></connection>
<connection>
<GID>210</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-62.5,145.5,-62.5</points>
<connection>
<GID>212</GID>
<name>IN_2</name></connection>
<connection>
<GID>210</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-63.5,145.5,-63.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<connection>
<GID>210</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-64.5,145.5,-64.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-55.5,148.5,-53.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<connection>
<GID>212</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153.5,-64.5,159.5,-64.5</points>
<connection>
<GID>228</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153.5,-63.5,159.5,-63.5</points>
<connection>
<GID>228</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>212</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-74.5,95.5,-49</points>
<connection>
<GID>209</GID>
<name>clock</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-74.5,148.5,-74.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>65.5 6</intersection>
<intersection>95.5 0</intersection>
<intersection>132.5 5</intersection>
<intersection>148.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>148.5,-74.5,148.5,-66.5</points>
<connection>
<GID>212</GID>
<name>clock</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>132.5,-74.5,132.5,-66.5</points>
<connection>
<GID>210</GID>
<name>clock</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>65.5,-74.5,65.5,-56</points>
<intersection>-74.5 1</intersection>
<intersection>-56 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>65.5,-56,71.5,-56</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>65.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-72.5,80.5,-49</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<connection>
<GID>208</GID>
<name>clear</name></connection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-72.5,150.5,-72.5</points>
<intersection>80.5 0</intersection>
<intersection>97.5 3</intersection>
<intersection>134.5 7</intersection>
<intersection>150.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-72.5,97.5,-49</points>
<connection>
<GID>209</GID>
<name>clear</name></connection>
<intersection>-72.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>150.5,-72.5,150.5,-66.5</points>
<connection>
<GID>212</GID>
<name>clear</name></connection>
<intersection>-72.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>134.5,-72.5,134.5,-66.5</points>
<connection>
<GID>210</GID>
<name>clear</name></connection>
<intersection>-72.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-41,119.5,-41</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>116.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-56,116.5,-41</points>
<connection>
<GID>211</GID>
<name>write_enable</name></connection>
<intersection>-56 4</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>104.5,-56,116.5,-56</points>
<connection>
<GID>234</GID>
<name>ENABLE_0</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-44,119.5,-44</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<connection>
<GID>211</GID>
<name>ENABLE_0</name></connection>
<intersection>119.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>119.5,-56,119.5,-44</points>
<intersection>-56 6</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>119.5,-56,125.5,-56</points>
<connection>
<GID>233</GID>
<name>ENABLE_0</name></connection>
<intersection>119.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-63.5,123.5,-63.5</points>
<connection>
<GID>234</GID>
<name>OUT_1</name></connection>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>114 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114,-63.5,114,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_1</name></connection>
<intersection>-63.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-62.5,123.5,-62.5</points>
<connection>
<GID>234</GID>
<name>OUT_2</name></connection>
<connection>
<GID>233</GID>
<name>IN_2</name></connection>
<intersection>113 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>113,-62.5,113,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_2</name></connection>
<intersection>-62.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-61.5,123.5,-61.5</points>
<connection>
<GID>234</GID>
<name>OUT_3</name></connection>
<connection>
<GID>233</GID>
<name>IN_3</name></connection>
<intersection>112 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>112,-61.5,112,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_3</name></connection>
<intersection>-61.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-60.5,123.5,-60.5</points>
<connection>
<GID>234</GID>
<name>OUT_4</name></connection>
<connection>
<GID>233</GID>
<name>IN_4</name></connection>
<intersection>111 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>111,-60.5,111,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_4</name></connection>
<intersection>-60.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-59.5,123.5,-59.5</points>
<connection>
<GID>234</GID>
<name>OUT_5</name></connection>
<connection>
<GID>233</GID>
<name>IN_5</name></connection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-59.5,110,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_5</name></connection>
<intersection>-59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-58.5,123.5,-58.5</points>
<connection>
<GID>234</GID>
<name>OUT_6</name></connection>
<connection>
<GID>233</GID>
<name>IN_6</name></connection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,-58.5,109,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_6</name></connection>
<intersection>-58.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-57.5,123.5,-57.5</points>
<connection>
<GID>234</GID>
<name>OUT_7</name></connection>
<connection>
<GID>233</GID>
<name>IN_7</name></connection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,-57.5,108,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_7</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-59.5,129.5,-59.5</points>
<connection>
<GID>233</GID>
<name>OUT_5</name></connection>
<connection>
<GID>210</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-64.5,129.5,-64.5</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-63.5,129.5,-63.5</points>
<connection>
<GID>233</GID>
<name>OUT_1</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-62.5,129.5,-62.5</points>
<connection>
<GID>233</GID>
<name>OUT_2</name></connection>
<connection>
<GID>210</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-61.5,129.5,-61.5</points>
<connection>
<GID>233</GID>
<name>OUT_3</name></connection>
<connection>
<GID>210</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-60.5,129.5,-60.5</points>
<connection>
<GID>233</GID>
<name>OUT_4</name></connection>
<connection>
<GID>210</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-57.5,129.5,-57.5</points>
<connection>
<GID>233</GID>
<name>OUT_7</name></connection>
<connection>
<GID>210</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-58.5,129.5,-58.5</points>
<connection>
<GID>233</GID>
<name>OUT_6</name></connection>
<connection>
<GID>210</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,-64.5,123.5,-64.5</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115,-64.5,115,-50.5</points>
<connection>
<GID>211</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>211</GID>
<name>DATA_IN_0</name></connection>
<intersection>-64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169.5,-61.5,171.5,-61.5</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<connection>
<GID>228</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-75.5,57,-75.5</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<connection>
<GID>215</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-73.5,57,-71.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-71.5,57,-71.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-57,78.5,-49</points>
<connection>
<GID>208</GID>
<name>clock</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-57,78.5,-57</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-58,71.5,-58</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>50.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50.5,-58,50.5,-55.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-38,78.5,-30</points>
<connection>
<GID>208</GID>
<name>load</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50.5,-49.5,50.5,-30</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-30,78.5,-30</points>
<intersection>50.5 1</intersection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-149,80,-147</points>
<intersection>-149 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-147,96.5,-147</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection>
<intersection>96.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-149,80,-149</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96.5,-147,96.5,-124</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-146,80,-123</points>
<intersection>-146 1</intersection>
<intersection>-125 2</intersection>
<intersection>-123 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-146,96.5,-146</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-125,80,-125</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-123,96.5,-123</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-147,80,-145</points>
<intersection>-147 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-145,96.5,-145</points>
<connection>
<GID>243</GID>
<name>IN_2</name></connection>
<intersection>80 0</intersection>
<intersection>96.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-147,80,-147</points>
<connection>
<GID>248</GID>
<name>OUT_1</name></connection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96.5,-145,96.5,-122</points>
<connection>
<GID>242</GID>
<name>IN_2</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-144,80,-121</points>
<intersection>-144 1</intersection>
<intersection>-123 2</intersection>
<intersection>-121 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-144,96.5,-144</points>
<connection>
<GID>243</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-123,80,-123</points>
<connection>
<GID>247</GID>
<name>OUT_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-121,96.5,-121</points>
<connection>
<GID>242</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-145,80,-143</points>
<intersection>-145 2</intersection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-143,96.5,-143</points>
<connection>
<GID>243</GID>
<name>IN_4</name></connection>
<intersection>80 0</intersection>
<intersection>96.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-145,80,-145</points>
<connection>
<GID>248</GID>
<name>OUT_2</name></connection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96.5,-143,96.5,-120</points>
<connection>
<GID>242</GID>
<name>IN_4</name></connection>
<intersection>-143 1</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-142,80,-119</points>
<intersection>-142 1</intersection>
<intersection>-121 2</intersection>
<intersection>-119 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-142,96.5,-142</points>
<connection>
<GID>243</GID>
<name>IN_5</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-121,80,-121</points>
<connection>
<GID>247</GID>
<name>OUT_2</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>80,-119,96.5,-119</points>
<connection>
<GID>242</GID>
<name>IN_5</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-143,80,-141</points>
<intersection>-143 2</intersection>
<intersection>-141 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-141,96.5,-141</points>
<connection>
<GID>243</GID>
<name>IN_6</name></connection>
<intersection>80 0</intersection>
<intersection>96.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-143,80,-143</points>
<connection>
<GID>248</GID>
<name>OUT_3</name></connection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96.5,-141,96.5,-118</points>
<connection>
<GID>242</GID>
<name>IN_6</name></connection>
<intersection>-141 1</intersection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-140,80,-117</points>
<intersection>-140 1</intersection>
<intersection>-119 2</intersection>
<intersection>-117 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-140,96.5,-140</points>
<connection>
<GID>243</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-119,80,-119</points>
<connection>
<GID>247</GID>
<name>OUT_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-117,96.5,-117</points>
<connection>
<GID>242</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-139,80,-116</points>
<intersection>-139 1</intersection>
<intersection>-137 2</intersection>
<intersection>-116 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-139,96.5,-139</points>
<connection>
<GID>243</GID>
<name>IN_8</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-137,80,-137</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>80,-116,96.5,-116</points>
<connection>
<GID>242</GID>
<name>IN_8</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-138,80,-113</points>
<intersection>-138 1</intersection>
<intersection>-115 4</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-138,96.5,-138</points>
<connection>
<GID>243</GID>
<name>IN_9</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-113,80,-113</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>80,-115,96.5,-115</points>
<connection>
<GID>242</GID>
<name>IN_9</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-137,80,-114</points>
<intersection>-137 1</intersection>
<intersection>-135 2</intersection>
<intersection>-114 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-137,96.5,-137</points>
<connection>
<GID>243</GID>
<name>IN_10</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-135,80,-135</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>80,-114,96.5,-114</points>
<connection>
<GID>242</GID>
<name>IN_10</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-136,80,-111</points>
<intersection>-136 1</intersection>
<intersection>-113 3</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-136,96.5,-136</points>
<connection>
<GID>243</GID>
<name>IN_11</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-111,80,-111</points>
<connection>
<GID>245</GID>
<name>OUT_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-113,96.5,-113</points>
<connection>
<GID>242</GID>
<name>IN_11</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-135,80,-112</points>
<intersection>-135 1</intersection>
<intersection>-133 2</intersection>
<intersection>-112 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-135,96.5,-135</points>
<connection>
<GID>243</GID>
<name>IN_12</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-133,80,-133</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-112,96.5,-112</points>
<connection>
<GID>242</GID>
<name>IN_12</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-134,80,-109</points>
<intersection>-134 1</intersection>
<intersection>-111 3</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-134,96.5,-134</points>
<connection>
<GID>243</GID>
<name>IN_13</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-109,80,-109</points>
<connection>
<GID>245</GID>
<name>OUT_2</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-111,96.5,-111</points>
<connection>
<GID>242</GID>
<name>IN_13</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-133,80,-110</points>
<intersection>-133 1</intersection>
<intersection>-131 2</intersection>
<intersection>-110 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-133,96.5,-133</points>
<connection>
<GID>243</GID>
<name>IN_14</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-131,80,-131</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-110,96.5,-110</points>
<connection>
<GID>242</GID>
<name>IN_14</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-132,80,-107</points>
<intersection>-132 1</intersection>
<intersection>-109 3</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-132,96.5,-132</points>
<connection>
<GID>243</GID>
<name>IN_15</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-107,80,-107</points>
<connection>
<GID>245</GID>
<name>OUT_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-109,96.5,-109</points>
<connection>
<GID>242</GID>
<name>IN_15</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-98.5,87,-98.5</points>
<connection>
<GID>253</GID>
<name>ENABLE</name></connection>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-93,138.5,-93</points>
<intersection>82.5 8</intersection>
<intersection>138.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>138.5,-144.5,138.5,-93</points>
<intersection>-144.5 18</intersection>
<intersection>-139.5 19</intersection>
<intersection>-134.5 20</intersection>
<intersection>-129.5 21</intersection>
<intersection>-124.5 22</intersection>
<intersection>-119.5 23</intersection>
<intersection>-114.5 24</intersection>
<intersection>-109.5 25</intersection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>82.5,-101.5,82.5,-93</points>
<intersection>-101.5 10</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>82.5,-101.5,87,-101.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>82.5 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>138.5,-144.5,141.5,-144.5</points>
<connection>
<GID>281</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>138.5,-139.5,141.5,-139.5</points>
<connection>
<GID>280</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>138.5,-134.5,141.5,-134.5</points>
<connection>
<GID>279</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>138.5,-129.5,141.5,-129.5</points>
<connection>
<GID>278</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>138.5,-124.5,141.5,-124.5</points>
<connection>
<GID>277</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>138.5,-119.5,141.5,-119.5</points>
<connection>
<GID>276</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>138.5,-114.5,141.5,-114.5</points>
<connection>
<GID>275</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>138.5,-109.5,141.5,-109.5</points>
<connection>
<GID>274</GID>
<name>SEL_0</name></connection>
<intersection>138.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-130.5,94,-101.5</points>
<intersection>-130.5 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-101.5,94,-101.5</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-130.5,98.5,-130.5</points>
<connection>
<GID>243</GID>
<name>ENABLE_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-107.5,98.5,-100.5</points>
<connection>
<GID>242</GID>
<name>ENABLE_0</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-100.5,98.5,-100.5</points>
<connection>
<GID>253</GID>
<name>OUT_1</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-143.5,115,-143.5</points>
<connection>
<GID>258</GID>
<name>carry_out</name></connection>
<connection>
<GID>259</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-147,102,-130.5</points>
<intersection>-147 2</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-130.5,112,-130.5</points>
<connection>
<GID>258</GID>
<name>IN_B_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-147,102,-147</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-145,102.5,-131.5</points>
<intersection>-145 2</intersection>
<intersection>-131.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-131.5,112,-131.5</points>
<connection>
<GID>258</GID>
<name>IN_B_1</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-145,102.5,-145</points>
<connection>
<GID>243</GID>
<name>OUT_2</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-143,103,-132.5</points>
<intersection>-143 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-132.5,112,-132.5</points>
<connection>
<GID>258</GID>
<name>IN_B_2</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-143,103,-143</points>
<connection>
<GID>243</GID>
<name>OUT_4</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-141,103.5,-133.5</points>
<intersection>-141 2</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-133.5,112,-133.5</points>
<connection>
<GID>258</GID>
<name>IN_B_3</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-141,103.5,-141</points>
<connection>
<GID>243</GID>
<name>OUT_6</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-146.5,105.5,-139</points>
<intersection>-146.5 1</intersection>
<intersection>-139 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-146.5,112,-146.5</points>
<connection>
<GID>259</GID>
<name>IN_B_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-139,105.5,-139</points>
<connection>
<GID>243</GID>
<name>OUT_8</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-147.5,105,-137</points>
<intersection>-147.5 1</intersection>
<intersection>-137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-147.5,112,-147.5</points>
<connection>
<GID>259</GID>
<name>IN_B_1</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-137,105,-137</points>
<connection>
<GID>243</GID>
<name>OUT_10</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-148.5,104.5,-135</points>
<intersection>-148.5 1</intersection>
<intersection>-135 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-148.5,112,-148.5</points>
<connection>
<GID>259</GID>
<name>IN_B_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-135,104.5,-135</points>
<connection>
<GID>243</GID>
<name>OUT_12</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-149.5,104,-133</points>
<intersection>-149.5 1</intersection>
<intersection>-133 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-149.5,112,-149.5</points>
<connection>
<GID>259</GID>
<name>IN_B_3</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-133,104,-133</points>
<connection>
<GID>243</GID>
<name>OUT_14</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-146,106,-137.5</points>
<intersection>-146 2</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-137.5,112,-137.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-146,106,-146</points>
<connection>
<GID>243</GID>
<name>OUT_1</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-144,106,-138.5</points>
<intersection>-144 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-138.5,112,-138.5</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-144,106,-144</points>
<connection>
<GID>243</GID>
<name>OUT_3</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-142,106,-139.5</points>
<intersection>-142 2</intersection>
<intersection>-139.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-139.5,112,-139.5</points>
<connection>
<GID>258</GID>
<name>IN_2</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-142,106,-142</points>
<connection>
<GID>243</GID>
<name>OUT_5</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-140.5,106,-140</points>
<intersection>-140.5 1</intersection>
<intersection>-140 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-140.5,112,-140.5</points>
<connection>
<GID>258</GID>
<name>IN_3</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-140,106,-140</points>
<connection>
<GID>243</GID>
<name>OUT_7</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-153.5,108,-138</points>
<intersection>-153.5 1</intersection>
<intersection>-138 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-153.5,112,-153.5</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-138,108,-138</points>
<connection>
<GID>243</GID>
<name>OUT_9</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-154.5,107.5,-136</points>
<intersection>-154.5 1</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-154.5,112,-154.5</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-136,107.5,-136</points>
<connection>
<GID>243</GID>
<name>OUT_11</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-155.5,107,-134</points>
<intersection>-155.5 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-155.5,112,-155.5</points>
<connection>
<GID>259</GID>
<name>IN_2</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-134,107,-134</points>
<connection>
<GID>243</GID>
<name>OUT_13</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-156.5,106.5,-132</points>
<intersection>-156.5 1</intersection>
<intersection>-132 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-156.5,112,-156.5</points>
<connection>
<GID>259</GID>
<name>IN_3</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-132,106.5,-132</points>
<connection>
<GID>243</GID>
<name>OUT_15</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-126,101.5,-124</points>
<intersection>-126 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-126,108.5,-126</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-124,101.5,-124</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-124,108.5,-124</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-124,100.5,-123</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>-124 1</intersection></vsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-122.5,104,-122</points>
<intersection>-122.5 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-122.5,113.5,-122.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-122,104,-122</points>
<connection>
<GID>242</GID>
<name>OUT_2</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-120.5,113.5,-120.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-121,100.5,-120.5</points>
<connection>
<GID>242</GID>
<name>OUT_3</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>100.5,-119,108.5,-119</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-120,100.5,-119</points>
<connection>
<GID>242</GID>
<name>OUT_4</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-119,101.5,-117</points>
<intersection>-119 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-117,108.5,-117</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-119,101.5,-119</points>
<connection>
<GID>242</GID>
<name>OUT_5</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-118,102.5,-115.5</points>
<intersection>-118 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,-115.5,113.5,-115.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-118,102.5,-118</points>
<connection>
<GID>242</GID>
<name>OUT_6</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-117,102,-113.5</points>
<intersection>-117 2</intersection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-113.5,113.5,-113.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-117,102,-117</points>
<connection>
<GID>242</GID>
<name>OUT_7</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-116,101.5,-112</points>
<intersection>-116 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-112,108.5,-112</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-116,101.5,-116</points>
<connection>
<GID>242</GID>
<name>OUT_8</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-115,101.5,-110</points>
<intersection>-115 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-110,108.5,-110</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-115,101.5,-115</points>
<connection>
<GID>242</GID>
<name>OUT_9</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-114,102,-108.5</points>
<intersection>-114 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-108.5,113.5,-108.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-114,102,-114</points>
<connection>
<GID>242</GID>
<name>OUT_10</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-113,102,-106.5</points>
<intersection>-113 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-106.5,113.5,-106.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-113,102,-113</points>
<connection>
<GID>242</GID>
<name>OUT_11</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-112,101.5,-105</points>
<intersection>-112 2</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-105,108.5,-105</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-112,101.5,-112</points>
<connection>
<GID>242</GID>
<name>OUT_12</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-111,101.5,-103</points>
<intersection>-111 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-103,108.5,-103</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-111,101.5,-111</points>
<connection>
<GID>242</GID>
<name>OUT_13</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-110,101,-101.5</points>
<intersection>-110 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-101.5,113.5,-101.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-110,101,-110</points>
<connection>
<GID>242</GID>
<name>OUT_14</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-109,100.5,-99.5</points>
<connection>
<GID>242</GID>
<name>OUT_15</name></connection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-99.5,113.5,-99.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-148,129.5,-134</points>
<intersection>-148 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-148,139.5,-148</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-134,129.5,-134</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-239.556,773.472,1538.44,-143.528</PageViewport>
<gate>
<ID>386</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-93</position>
<output>
<ID>OUT_0</ID>545 </output>
<output>
<ID>OUT_1</ID>547 </output>
<output>
<ID>OUT_2</ID>549 </output>
<output>
<ID>OUT_3</ID>551 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>387</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-117</position>
<output>
<ID>OUT_0</ID>544 </output>
<output>
<ID>OUT_1</ID>546 </output>
<output>
<ID>OUT_2</ID>548 </output>
<output>
<ID>OUT_3</ID>550 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>-35.5,-106</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>389</ID>
<type>AA_LABEL</type>
<position>-36,-80</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>AA_LABEL</type>
<position>-36,-92.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>AA_LABEL</type>
<position>-36,-117.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>BA_DECODER_2x4</type>
<position>5.5,-71</position>
<input>
<ID>ENABLE</ID>560 </input>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>562 </output>
<output>
<ID>OUT_1</ID>563 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_TOGGLE</type>
<position>0.5,-69.5</position>
<output>
<ID>OUT_0</ID>560 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_TOGGLE</type>
<position>-4,-72.5</position>
<output>
<ID>OUT_0</ID>561 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_LABEL</type>
<position>1,-66.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_LABEL</type>
<position>-10.5,-72</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,-106.5</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>574 </input>
<input>
<ID>IN_2</ID>575 </input>
<input>
<ID>IN_3</ID>576 </input>
<input>
<ID>IN_B_0</ID>565 </input>
<input>
<ID>IN_B_1</ID>566 </input>
<input>
<ID>IN_B_2</ID>567 </input>
<input>
<ID>IN_B_3</ID>568 </input>
<output>
<ID>OUT_0</ID>597 </output>
<output>
<ID>OUT_1</ID>598 </output>
<output>
<ID>OUT_2</ID>599 </output>
<output>
<ID>OUT_3</ID>600 </output>
<output>
<ID>carry_out</ID>564 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>398</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,-122.5</position>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>578 </input>
<input>
<ID>IN_2</ID>579 </input>
<input>
<ID>IN_3</ID>580 </input>
<input>
<ID>IN_B_0</ID>569 </input>
<input>
<ID>IN_B_1</ID>570 </input>
<input>
<ID>IN_B_2</ID>571 </input>
<input>
<ID>IN_B_3</ID>572 </input>
<output>
<ID>OUT_0</ID>601 </output>
<output>
<ID>OUT_1</ID>602 </output>
<output>
<ID>OUT_2</ID>603 </output>
<output>
<ID>OUT_3</ID>604 </output>
<input>
<ID>carry_in</ID>564 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>399</ID>
<type>AA_LABEL</type>
<position>39,-99</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>39.5,-127.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_LABEL</type>
<position>25,-100</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>AA_LABEL</type>
<position>25.5,-106.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AA_LABEL</type>
<position>25,-116</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>AA_LABEL</type>
<position>26,-123</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>27,-96</position>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>32,-92.5</position>
<input>
<ID>IN_0</ID>584 </input>
<input>
<ID>IN_1</ID>583 </input>
<output>
<ID>OUT</ID>606 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>27,-89</position>
<input>
<ID>IN_0</ID>586 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>32,-85.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>587 </input>
<output>
<ID>OUT</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>27,-82</position>
<input>
<ID>IN_0</ID>590 </input>
<input>
<ID>IN_1</ID>589 </input>
<output>
<ID>OUT</ID>609 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>32,-78.5</position>
<input>
<ID>IN_0</ID>592 </input>
<input>
<ID>IN_1</ID>591 </input>
<output>
<ID>OUT</ID>610 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_AND2</type>
<position>27,-75</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>593 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_AND2</type>
<position>32,-71.5</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>595 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>413</ID>
<type>AA_MUX_2x1</type>
<position>57,-83</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>612 </input>
<output>
<ID>OUT</ID>620 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>AA_MUX_2x1</type>
<position>57,-88</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>611 </input>
<output>
<ID>OUT</ID>619 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_MUX_2x1</type>
<position>57,-93</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>610 </input>
<output>
<ID>OUT</ID>618 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_MUX_2x1</type>
<position>57,-98</position>
<input>
<ID>IN_0</ID>601 </input>
<input>
<ID>IN_1</ID>609 </input>
<output>
<ID>OUT</ID>617 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>AA_MUX_2x1</type>
<position>57,-103</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>608 </input>
<output>
<ID>OUT</ID>616 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_MUX_2x1</type>
<position>57,-108</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>615 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_MUX_2x1</type>
<position>57,-113</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>614 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_MUX_2x1</type>
<position>57,-118</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>605 </input>
<output>
<ID>OUT</ID>613 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>79.5,-100</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>614 </input>
<input>
<ID>IN_2</ID>615 </input>
<input>
<ID>IN_3</ID>616 </input>
<input>
<ID>IN_4</ID>617 </input>
<input>
<ID>IN_5</ID>618 </input>
<input>
<ID>IN_6</ID>619 </input>
<input>
<ID>IN_7</ID>620 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 54</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>422</ID>
<type>AA_LABEL</type>
<position>57,-121.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>58,-79</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>424</ID>
<type>GA_LED</type>
<position>71,-110</position>
<input>
<ID>N_in2</ID>620 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>425</ID>
<type>GA_LED</type>
<position>73.5,-110</position>
<input>
<ID>N_in2</ID>619 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>426</ID>
<type>GA_LED</type>
<position>76,-110</position>
<input>
<ID>N_in2</ID>618 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>427</ID>
<type>GA_LED</type>
<position>78.5,-110</position>
<input>
<ID>N_in2</ID>617 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>428</ID>
<type>GA_LED</type>
<position>81,-110</position>
<input>
<ID>N_in2</ID>616 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>429</ID>
<type>GA_LED</type>
<position>83.5,-110</position>
<input>
<ID>N_in2</ID>615 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>430</ID>
<type>GA_LED</type>
<position>86,-110</position>
<input>
<ID>N_in2</ID>614 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>431</ID>
<type>GA_LED</type>
<position>88.5,-110</position>
<input>
<ID>N_in2</ID>613 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>88.5,-112</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AA_LABEL</type>
<position>86,-112</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>83.5,-112</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>81,-112</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>78.5,-112</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AA_LABEL</type>
<position>76,-112</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>73.5,-112</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>71,-112</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>207,-63.5</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>AA_LABEL</type>
<position>207,-74.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>AE_REGISTER8</type>
<position>150,-74.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>644 </output>
<output>
<ID>OUT_1</ID>643 </output>
<output>
<ID>OUT_2</ID>642 </output>
<output>
<ID>OUT_3</ID>641 </output>
<output>
<ID>OUT_4</ID>640 </output>
<output>
<ID>OUT_5</ID>639 </output>
<output>
<ID>OUT_6</ID>638 </output>
<output>
<ID>OUT_7</ID>637 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>684 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>443</ID>
<type>AE_REGISTER8</type>
<position>150,-87.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>660 </output>
<output>
<ID>OUT_1</ID>651 </output>
<output>
<ID>OUT_2</ID>650 </output>
<output>
<ID>OUT_3</ID>649 </output>
<output>
<ID>OUT_4</ID>648 </output>
<output>
<ID>OUT_5</ID>647 </output>
<output>
<ID>OUT_6</ID>646 </output>
<output>
<ID>OUT_7</ID>645 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>685 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>444</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-37</position>
<input>
<ID>IN_0</ID>645 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>621 </input>
<output>
<ID>OUT</ID>652 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>445</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-48</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>638 </input>
<input>
<ID>IN_2</ID>630 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>653 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>446</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-59</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>639 </input>
<input>
<ID>IN_2</ID>631 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT</ID>654 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>447</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-68.5</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>640 </input>
<input>
<ID>IN_2</ID>632 </input>
<input>
<ID>IN_3</ID>624 </input>
<output>
<ID>OUT</ID>655 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-79.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>641 </input>
<input>
<ID>IN_2</ID>633 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT</ID>656 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-90.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>642 </input>
<input>
<ID>IN_2</ID>634 </input>
<input>
<ID>IN_3</ID>626 </input>
<output>
<ID>OUT</ID>657 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>450</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-101</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>643 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>658 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>451</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-112</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>644 </input>
<input>
<ID>IN_2</ID>636 </input>
<input>
<ID>IN_3</ID>628 </input>
<output>
<ID>OUT</ID>659 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>452</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>207.5,-69.5</position>
<input>
<ID>IN_0</ID>659 </input>
<input>
<ID>IN_1</ID>658 </input>
<input>
<ID>IN_2</ID>657 </input>
<input>
<ID>IN_3</ID>656 </input>
<input>
<ID>IN_4</ID>655 </input>
<input>
<ID>IN_5</ID>654 </input>
<input>
<ID>IN_6</ID>653 </input>
<input>
<ID>IN_7</ID>652 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>453</ID>
<type>DD_KEYPAD_HEX</type>
<position>117,-52</position>
<output>
<ID>OUT_0</ID>662 </output>
<output>
<ID>OUT_1</ID>663 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>454</ID>
<type>BB_CLOCK</type>
<position>138.5,-96</position>
<output>
<ID>CLK</ID>661 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>151,-41</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>151,-54</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_LABEL</type>
<position>151,-67.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AA_LABEL</type>
<position>151,-80.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>459</ID>
<type>AA_LABEL</type>
<position>115.5,-45</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>460</ID>
<type>DD_KEYPAD_HEX</type>
<position>117,-66</position>
<output>
<ID>OUT_0</ID>672 </output>
<output>
<ID>OUT_1</ID>673 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_MUX_4x1</type>
<position>188,-37</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>621 </input>
<output>
<ID>OUT</ID>664 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_MUX_4x1</type>
<position>188,-48</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>638 </input>
<input>
<ID>IN_2</ID>630 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>665 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_MUX_4x1</type>
<position>188,-59</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>639 </input>
<input>
<ID>IN_2</ID>631 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT</ID>666 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_MUX_4x1</type>
<position>188,-68.5</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>640 </input>
<input>
<ID>IN_2</ID>632 </input>
<input>
<ID>IN_3</ID>624 </input>
<output>
<ID>OUT</ID>667 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>465</ID>
<type>AE_MUX_4x1</type>
<position>188,-79.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>641 </input>
<input>
<ID>IN_2</ID>633 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT</ID>668 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>466</ID>
<type>AE_MUX_4x1</type>
<position>188,-90.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>642 </input>
<input>
<ID>IN_2</ID>634 </input>
<input>
<ID>IN_3</ID>626 </input>
<output>
<ID>OUT</ID>669 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_MUX_4x1</type>
<position>188,-101</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>643 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>670 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>468</ID>
<type>AE_MUX_4x1</type>
<position>188,-112</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>644 </input>
<input>
<ID>IN_2</ID>636 </input>
<input>
<ID>IN_3</ID>628 </input>
<output>
<ID>OUT</ID>671 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>469</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>207.5,-80.5</position>
<input>
<ID>IN_0</ID>671 </input>
<input>
<ID>IN_1</ID>670 </input>
<input>
<ID>IN_2</ID>669 </input>
<input>
<ID>IN_3</ID>668 </input>
<input>
<ID>IN_4</ID>667 </input>
<input>
<ID>IN_5</ID>666 </input>
<input>
<ID>IN_6</ID>665 </input>
<input>
<ID>IN_7</ID>664 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_LABEL</type>
<position>115.5,-59</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>DD_KEYPAD_HEX</type>
<position>133,-65.5</position>
<output>
<ID>OUT_0</ID>677 </output>
<output>
<ID>OUT_1</ID>676 </output>
<output>
<ID>OUT_2</ID>675 </output>
<output>
<ID>OUT_3</ID>674 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>472</ID>
<type>DD_KEYPAD_HEX</type>
<position>133,-77.5</position>
<output>
<ID>OUT_0</ID>681 </output>
<output>
<ID>OUT_1</ID>680 </output>
<output>
<ID>OUT_2</ID>679 </output>
<output>
<ID>OUT_3</ID>678 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>473</ID>
<type>AA_LABEL</type>
<position>133,-58.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>BA_DECODER_2x4</type>
<position>135,-32.5</position>
<input>
<ID>ENABLE</ID>686 </input>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>688 </input>
<output>
<ID>OUT_0</ID>682 </output>
<output>
<ID>OUT_1</ID>683 </output>
<output>
<ID>OUT_2</ID>684 </output>
<output>
<ID>OUT_3</ID>685 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_TOGGLE</type>
<position>129,-32</position>
<output>
<ID>OUT_0</ID>686 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>476</ID>
<type>AA_LABEL</type>
<position>126.5,-30.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>477</ID>
<type>DD_KEYPAD_HEX</type>
<position>130,-45</position>
<output>
<ID>OUT_0</ID>687 </output>
<output>
<ID>OUT_1</ID>688 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>130.5,-38</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>AE_REGISTER8</type>
<position>150,-48</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>628 </output>
<output>
<ID>OUT_1</ID>627 </output>
<output>
<ID>OUT_2</ID>626 </output>
<output>
<ID>OUT_3</ID>625 </output>
<output>
<ID>OUT_4</ID>624 </output>
<output>
<ID>OUT_5</ID>623 </output>
<output>
<ID>OUT_6</ID>622 </output>
<output>
<ID>OUT_7</ID>621 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>682 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>480</ID>
<type>AE_REGISTER8</type>
<position>150,-61</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>636 </output>
<output>
<ID>OUT_1</ID>635 </output>
<output>
<ID>OUT_2</ID>634 </output>
<output>
<ID>OUT_3</ID>633 </output>
<output>
<ID>OUT_4</ID>632 </output>
<output>
<ID>OUT_5</ID>631 </output>
<output>
<ID>OUT_6</ID>630 </output>
<output>
<ID>OUT_7</ID>629 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>683 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>481</ID>
<type>AA_LABEL</type>
<position>160.5,-23.5</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>483</ID>
<type>AA_LABEL</type>
<position>19.5,-37</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>485</ID>
<type>AA_LABEL</type>
<position>96,37.5</position>
<gparam>LABEL_TEXT Last update before starting to connect the pieces</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>87.5,20.5</position>
<gparam>LABEL_TEXT Check page 6</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>AA_INVERTER</type>
<position>-34,-23.5</position>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>543 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_TOGGLE</type>
<position>-9.5,1</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_LABEL</type>
<position>-32,-31</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>AA_LABEL</type>
<position>-32,-32.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AE_REGISTER8</type>
<position>-5,-15</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>481 </input>
<input>
<ID>IN_2</ID>482 </input>
<input>
<ID>IN_3</ID>483 </input>
<input>
<ID>IN_4</ID>484 </input>
<input>
<ID>IN_5</ID>485 </input>
<input>
<ID>IN_6</ID>486 </input>
<input>
<ID>IN_7</ID>487 </input>
<output>
<ID>OUT_0</ID>495 </output>
<output>
<ID>OUT_1</ID>494 </output>
<output>
<ID>OUT_2</ID>493 </output>
<output>
<ID>OUT_3</ID>492 </output>
<output>
<ID>OUT_4</ID>491 </output>
<output>
<ID>OUT_5</ID>490 </output>
<output>
<ID>OUT_6</ID>489 </output>
<output>
<ID>OUT_7</ID>488 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>541 </input>
<input>
<ID>count_enable</ID>503 </input>
<input>
<ID>count_up</ID>503 </input>
<input>
<ID>load</ID>543 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>348</ID>
<type>AE_REGISTER8</type>
<position>12,-15</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>494 </input>
<input>
<ID>IN_2</ID>493 </input>
<input>
<ID>IN_3</ID>492 </input>
<input>
<ID>IN_4</ID>491 </input>
<input>
<ID>IN_5</ID>490 </input>
<input>
<ID>IN_6</ID>489 </input>
<input>
<ID>IN_7</ID>488 </input>
<output>
<ID>OUT_0</ID>506 </output>
<output>
<ID>OUT_1</ID>505 </output>
<output>
<ID>OUT_2</ID>501 </output>
<output>
<ID>OUT_3</ID>500 </output>
<output>
<ID>OUT_4</ID>499 </output>
<output>
<ID>OUT_5</ID>498 </output>
<output>
<ID>OUT_6</ID>497 </output>
<output>
<ID>OUT_7</ID>496 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>502 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>349</ID>
<type>AE_REGISTER8</type>
<position>49,-32.5</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>531 </input>
<input>
<ID>IN_2</ID>532 </input>
<input>
<ID>IN_3</ID>533 </input>
<input>
<ID>IN_4</ID>534 </input>
<input>
<ID>IN_5</ID>529 </input>
<input>
<ID>IN_6</ID>536 </input>
<input>
<ID>IN_7</ID>535 </input>
<output>
<ID>OUT_0</ID>514 </output>
<output>
<ID>OUT_1</ID>513 </output>
<output>
<ID>OUT_2</ID>512 </output>
<output>
<ID>OUT_3</ID>511 </output>
<output>
<ID>OUT_4</ID>510 </output>
<output>
<ID>OUT_5</ID>509 </output>
<output>
<ID>OUT_6</ID>508 </output>
<output>
<ID>OUT_7</ID>507 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>504 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_RAM_8x8</type>
<position>27,-14.5</position>
<input>
<ID>ADDRESS_0</ID>506 </input>
<input>
<ID>ADDRESS_1</ID>505 </input>
<input>
<ID>ADDRESS_2</ID>501 </input>
<input>
<ID>ADDRESS_3</ID>500 </input>
<input>
<ID>ADDRESS_4</ID>499 </input>
<input>
<ID>ADDRESS_5</ID>498 </input>
<input>
<ID>ADDRESS_6</ID>497 </input>
<input>
<ID>ADDRESS_7</ID>496 </input>
<input>
<ID>DATA_IN_0</ID>537 </input>
<input>
<ID>DATA_IN_1</ID>522 </input>
<input>
<ID>DATA_IN_2</ID>523 </input>
<input>
<ID>DATA_IN_3</ID>524 </input>
<input>
<ID>DATA_IN_4</ID>525 </input>
<input>
<ID>DATA_IN_5</ID>526 </input>
<input>
<ID>DATA_IN_6</ID>527 </input>
<input>
<ID>DATA_IN_7</ID>528 </input>
<output>
<ID>DATA_OUT_0</ID>537 </output>
<output>
<ID>DATA_OUT_1</ID>522 </output>
<output>
<ID>DATA_OUT_2</ID>523 </output>
<output>
<ID>DATA_OUT_3</ID>524 </output>
<output>
<ID>DATA_OUT_4</ID>525 </output>
<output>
<ID>DATA_OUT_5</ID>526 </output>
<output>
<ID>DATA_OUT_6</ID>527 </output>
<output>
<ID>DATA_OUT_7</ID>528 </output>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>write_enable</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_REGISTER8</type>
<position>65,-32.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>513 </input>
<input>
<ID>IN_2</ID>512 </input>
<input>
<ID>IN_3</ID>511 </input>
<input>
<ID>IN_4</ID>510 </input>
<input>
<ID>IN_5</ID>509 </input>
<input>
<ID>IN_6</ID>508 </input>
<input>
<ID>IN_7</ID>507 </input>
<output>
<ID>OUT_0</ID>516 </output>
<output>
<ID>OUT_1</ID>517 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>515 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>352</ID>
<type>DD_KEYPAD_HEX</type>
<position>-24.5,-21</position>
<output>
<ID>OUT_0</ID>480 </output>
<output>
<ID>OUT_1</ID>481 </output>
<output>
<ID>OUT_2</ID>482 </output>
<output>
<ID>OUT_3</ID>483 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>353</ID>
<type>DD_KEYPAD_HEX</type>
<position>-24.5,-9</position>
<output>
<ID>OUT_0</ID>484 </output>
<output>
<ID>OUT_1</ID>485 </output>
<output>
<ID>OUT_2</ID>486 </output>
<output>
<ID>OUT_3</ID>487 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>354</ID>
<type>BB_CLOCK</type>
<position>-36,-46.5</position>
<output>
<ID>CLK</ID>539 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_TOGGLE</type>
<position>-7,4</position>
<output>
<ID>OUT_0</ID>503 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>-19.5,2</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>357</ID>
<type>AA_LABEL</type>
<position>-19.5,4.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>6,1.5</position>
<output>
<ID>OUT_0</ID>502 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_TOGGLE</type>
<position>-6,-43.5</position>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_LABEL</type>
<position>-11.5,-40.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>AA_TOGGLE</type>
<position>45,-25</position>
<output>
<ID>OUT_0</ID>504 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>-10,-7</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>6.5,-7</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>27,-6</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>49,-22</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_TOGGLE</type>
<position>62,-24.5</position>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>367</ID>
<type>BE_ROM_8x8</type>
<position>80,-32</position>
<input>
<ID>ADDRESS_0</ID>516 </input>
<input>
<ID>ADDRESS_1</ID>517 </input>
<input>
<ID>ENABLE_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>368</ID>
<type>AA_TOGGLE</type>
<position>37,-12</position>
<output>
<ID>OUT_0</ID>520 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_TOGGLE</type>
<position>37,-15</position>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>43.5,-11.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>AA_LABEL</type>
<position>44,-14.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>41,-32</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>522 </input>
<input>
<ID>IN_2</ID>523 </input>
<input>
<ID>IN_3</ID>524 </input>
<input>
<ID>IN_4</ID>525 </input>
<input>
<ID>IN_5</ID>526 </input>
<input>
<ID>IN_6</ID>527 </input>
<input>
<ID>IN_7</ID>528 </input>
<output>
<ID>OUT_0</ID>530 </output>
<output>
<ID>OUT_1</ID>531 </output>
<output>
<ID>OUT_2</ID>532 </output>
<output>
<ID>OUT_3</ID>533 </output>
<output>
<ID>OUT_4</ID>534 </output>
<output>
<ID>OUT_5</ID>529 </output>
<output>
<ID>OUT_6</ID>536 </output>
<output>
<ID>OUT_7</ID>535 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>373</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>20,-32</position>
<input>
<ID>ENABLE_0</ID>520 </input>
<output>
<ID>OUT_0</ID>537 </output>
<output>
<ID>OUT_1</ID>522 </output>
<output>
<ID>OUT_2</ID>523 </output>
<output>
<ID>OUT_3</ID>524 </output>
<output>
<ID>OUT_4</ID>525 </output>
<output>
<ID>OUT_5</ID>526 </output>
<output>
<ID>OUT_6</ID>527 </output>
<output>
<ID>OUT_7</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_LABEL</type>
<position>66.5,-24</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>375</ID>
<type>AA_TOGGLE</type>
<position>89,-32.5</position>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>376</ID>
<type>AA_LABEL</type>
<position>90.5,-29.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND2</type>
<position>-10,-28</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>542 </input>
<output>
<ID>OUT</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_AND2</type>
<position>-24.5,-45.5</position>
<input>
<ID>IN_0</ID>540 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AA_TOGGLE</type>
<position>-30,-42.5</position>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_TOGGLE</type>
<position>-39,-29</position>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>381</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>14,-87.5</position>
<input>
<ID>ENABLE_0</ID>563 </input>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>545 </input>
<input>
<ID>IN_10</ID>554 </input>
<input>
<ID>IN_11</ID>555 </input>
<input>
<ID>IN_12</ID>556 </input>
<input>
<ID>IN_13</ID>557 </input>
<input>
<ID>IN_14</ID>558 </input>
<input>
<ID>IN_15</ID>559 </input>
<input>
<ID>IN_2</ID>546 </input>
<input>
<ID>IN_3</ID>547 </input>
<input>
<ID>IN_4</ID>548 </input>
<input>
<ID>IN_5</ID>549 </input>
<input>
<ID>IN_6</ID>550 </input>
<input>
<ID>IN_7</ID>551 </input>
<input>
<ID>IN_8</ID>552 </input>
<input>
<ID>IN_9</ID>553 </input>
<output>
<ID>OUT_0</ID>581 </output>
<output>
<ID>OUT_1</ID>582 </output>
<output>
<ID>OUT_10</ID>591 </output>
<output>
<ID>OUT_11</ID>592 </output>
<output>
<ID>OUT_12</ID>593 </output>
<output>
<ID>OUT_13</ID>594 </output>
<output>
<ID>OUT_14</ID>595 </output>
<output>
<ID>OUT_15</ID>596 </output>
<output>
<ID>OUT_2</ID>583 </output>
<output>
<ID>OUT_3</ID>584 </output>
<output>
<ID>OUT_4</ID>585 </output>
<output>
<ID>OUT_5</ID>586 </output>
<output>
<ID>OUT_6</ID>587 </output>
<output>
<ID>OUT_7</ID>588 </output>
<output>
<ID>OUT_8</ID>589 </output>
<output>
<ID>OUT_9</ID>590 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>382</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>14,-110.5</position>
<input>
<ID>ENABLE_0</ID>562 </input>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>545 </input>
<input>
<ID>IN_10</ID>554 </input>
<input>
<ID>IN_11</ID>555 </input>
<input>
<ID>IN_12</ID>556 </input>
<input>
<ID>IN_13</ID>557 </input>
<input>
<ID>IN_14</ID>558 </input>
<input>
<ID>IN_15</ID>559 </input>
<input>
<ID>IN_2</ID>546 </input>
<input>
<ID>IN_3</ID>547 </input>
<input>
<ID>IN_4</ID>548 </input>
<input>
<ID>IN_5</ID>549 </input>
<input>
<ID>IN_6</ID>550 </input>
<input>
<ID>IN_7</ID>551 </input>
<input>
<ID>IN_8</ID>552 </input>
<input>
<ID>IN_9</ID>553 </input>
<output>
<ID>OUT_0</ID>565 </output>
<output>
<ID>OUT_1</ID>573 </output>
<output>
<ID>OUT_10</ID>570 </output>
<output>
<ID>OUT_11</ID>578 </output>
<output>
<ID>OUT_12</ID>571 </output>
<output>
<ID>OUT_13</ID>579 </output>
<output>
<ID>OUT_14</ID>572 </output>
<output>
<ID>OUT_15</ID>580 </output>
<output>
<ID>OUT_2</ID>566 </output>
<output>
<ID>OUT_3</ID>574 </output>
<output>
<ID>OUT_4</ID>567 </output>
<output>
<ID>OUT_5</ID>575 </output>
<output>
<ID>OUT_6</ID>568 </output>
<output>
<ID>OUT_7</ID>576 </output>
<output>
<ID>OUT_8</ID>569 </output>
<output>
<ID>OUT_9</ID>577 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_LABEL</type>
<position>-8.5,-74.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-81</position>
<output>
<ID>OUT_0</ID>553 </output>
<output>
<ID>OUT_1</ID>555 </output>
<output>
<ID>OUT_2</ID>557 </output>
<output>
<ID>OUT_3</ID>559 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>385</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-105</position>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>554 </output>
<output>
<ID>OUT_2</ID>556 </output>
<output>
<ID>OUT_3</ID>558 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-24,-14.5,-18</points>
<intersection>-24 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-18,-9,-18</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-24,-14.5,-24</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-22,-14.5,-17</points>
<intersection>-22 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-17,-9,-17</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-22,-14.5,-22</points>
<connection>
<GID>352</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-20,-14.5,-16</points>
<intersection>-20 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-16,-9,-16</points>
<connection>
<GID>347</GID>
<name>IN_2</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-20,-14.5,-20</points>
<connection>
<GID>352</GID>
<name>OUT_2</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-18,-14.5,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-15,-9,-15</points>
<connection>
<GID>347</GID>
<name>IN_3</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-18,-14.5,-18</points>
<connection>
<GID>352</GID>
<name>OUT_3</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-14,-14.5,-12</points>
<intersection>-14 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-14,-9,-14</points>
<connection>
<GID>347</GID>
<name>IN_4</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-12,-14.5,-12</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-13,-14.5,-10</points>
<intersection>-13 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-13,-9,-13</points>
<connection>
<GID>347</GID>
<name>IN_5</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-10,-14.5,-10</points>
<connection>
<GID>353</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-12,-14.5,-8</points>
<intersection>-12 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-12,-9,-12</points>
<connection>
<GID>347</GID>
<name>IN_6</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-8,-14.5,-8</points>
<connection>
<GID>353</GID>
<name>OUT_2</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-11,-9,-11</points>
<connection>
<GID>347</GID>
<name>IN_7</name></connection>
<intersection>-19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19.5,-11,-19.5,-6</points>
<connection>
<GID>353</GID>
<name>OUT_3</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-11,8,-11</points>
<connection>
<GID>348</GID>
<name>IN_7</name></connection>
<connection>
<GID>347</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-12,8,-12</points>
<connection>
<GID>348</GID>
<name>IN_6</name></connection>
<connection>
<GID>347</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-13,8,-13</points>
<connection>
<GID>348</GID>
<name>IN_5</name></connection>
<connection>
<GID>347</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-14,8,-14</points>
<connection>
<GID>348</GID>
<name>IN_4</name></connection>
<connection>
<GID>347</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-15,8,-15</points>
<connection>
<GID>348</GID>
<name>IN_3</name></connection>
<connection>
<GID>347</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-16,8,-16</points>
<connection>
<GID>348</GID>
<name>IN_2</name></connection>
<connection>
<GID>347</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-17,8,-17</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<connection>
<GID>347</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-18,8,-18</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-11,22,-11</points>
<connection>
<GID>350</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>348</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-12,22,-12</points>
<connection>
<GID>350</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>348</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-13,22,-13</points>
<connection>
<GID>350</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>348</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-14,22,-14</points>
<connection>
<GID>350</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>348</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-15,22,-15</points>
<connection>
<GID>350</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>348</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-16,22,-16</points>
<connection>
<GID>350</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>348</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-9,11,1.5</points>
<connection>
<GID>348</GID>
<name>load</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,1.5,11,1.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-9,-5,4</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<connection>
<GID>347</GID>
<name>count_enable</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5,-8,-4,-8</points>
<intersection>-5 0</intersection>
<intersection>-4 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4,-9,-4,-8</points>
<connection>
<GID>347</GID>
<name>count_up</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>47,-25,48,-25</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-26.5,48,-25</points>
<connection>
<GID>349</GID>
<name>load</name></connection>
<intersection>-25 2</intersection></vsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-17,22,-17</points>
<connection>
<GID>350</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>348</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-18,22,-18</points>
<connection>
<GID>350</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-28.5,61,-28.5</points>
<connection>
<GID>351</GID>
<name>IN_7</name></connection>
<connection>
<GID>349</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-29.5,61,-29.5</points>
<connection>
<GID>351</GID>
<name>IN_6</name></connection>
<connection>
<GID>349</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-30.5,61,-30.5</points>
<connection>
<GID>351</GID>
<name>IN_5</name></connection>
<connection>
<GID>349</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-31.5,61,-31.5</points>
<connection>
<GID>351</GID>
<name>IN_4</name></connection>
<connection>
<GID>349</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-32.5,61,-32.5</points>
<connection>
<GID>351</GID>
<name>IN_3</name></connection>
<connection>
<GID>349</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-33.5,61,-33.5</points>
<connection>
<GID>351</GID>
<name>IN_2</name></connection>
<connection>
<GID>349</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-34.5,61,-34.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<connection>
<GID>349</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-35.5,61,-35.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-26.5,64,-24.5</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<connection>
<GID>351</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-35.5,75,-35.5</points>
<connection>
<GID>367</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-34.5,75,-34.5</points>
<connection>
<GID>367</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>351</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-45.5,11,-20</points>
<connection>
<GID>348</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-45.5,64,-45.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>-19 6</intersection>
<intersection>11 0</intersection>
<intersection>48 5</intersection>
<intersection>64 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>64,-45.5,64,-37.5</points>
<connection>
<GID>351</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>48,-45.5,48,-37.5</points>
<connection>
<GID>349</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-19,-45.5,-19,-27</points>
<intersection>-45.5 1</intersection>
<intersection>-27 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-19,-27,-13,-27</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-19 6</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-43.5,-4,-20</points>
<connection>
<GID>359</GID>
<name>OUT_0</name></connection>
<connection>
<GID>347</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4,-43.5,66,-43.5</points>
<intersection>-4 0</intersection>
<intersection>13 3</intersection>
<intersection>50 7</intersection>
<intersection>66 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-43.5,13,-20</points>
<connection>
<GID>348</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>66,-43.5,66,-37.5</points>
<connection>
<GID>351</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>50,-43.5,50,-37.5</points>
<connection>
<GID>349</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-12,35,-12</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-27,33,-12</points>
<intersection>-27 4</intersection>
<intersection>-14 7</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-27,33,-27</points>
<connection>
<GID>373</GID>
<name>ENABLE_0</name></connection>
<intersection>33 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>32,-14,33,-14</points>
<connection>
<GID>350</GID>
<name>write_enable</name></connection>
<intersection>33 3</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-15,35,-15</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>ENABLE_0</name></connection>
<intersection>35 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35,-27,35,-15</points>
<intersection>-27 6</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35,-27,41,-27</points>
<connection>
<GID>372</GID>
<name>ENABLE_0</name></connection>
<intersection>35 5</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-34.5,39,-34.5</points>
<connection>
<GID>373</GID>
<name>OUT_1</name></connection>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29.5,-34.5,29.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_1</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-33.5,39,-33.5</points>
<connection>
<GID>373</GID>
<name>OUT_2</name></connection>
<connection>
<GID>372</GID>
<name>IN_2</name></connection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-33.5,28.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_2</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-32.5,39,-32.5</points>
<connection>
<GID>373</GID>
<name>OUT_3</name></connection>
<connection>
<GID>372</GID>
<name>IN_3</name></connection>
<intersection>27.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>27.5,-32.5,27.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_3</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-31.5,39,-31.5</points>
<connection>
<GID>373</GID>
<name>OUT_4</name></connection>
<connection>
<GID>372</GID>
<name>IN_4</name></connection>
<intersection>26.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26.5,-31.5,26.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_4</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-30.5,39,-30.5</points>
<connection>
<GID>373</GID>
<name>OUT_5</name></connection>
<connection>
<GID>372</GID>
<name>IN_5</name></connection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-30.5,25.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_5</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-29.5,39,-29.5</points>
<connection>
<GID>373</GID>
<name>OUT_6</name></connection>
<connection>
<GID>372</GID>
<name>IN_6</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-29.5,24.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_6</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-28.5,39,-28.5</points>
<connection>
<GID>373</GID>
<name>OUT_7</name></connection>
<connection>
<GID>372</GID>
<name>IN_7</name></connection>
<intersection>23.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-28.5,23.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_7</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-30.5,45,-30.5</points>
<connection>
<GID>372</GID>
<name>OUT_5</name></connection>
<connection>
<GID>349</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-35.5,45,-35.5</points>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-34.5,45,-34.5</points>
<connection>
<GID>372</GID>
<name>OUT_1</name></connection>
<connection>
<GID>349</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-33.5,45,-33.5</points>
<connection>
<GID>372</GID>
<name>OUT_2</name></connection>
<connection>
<GID>349</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-32.5,45,-32.5</points>
<connection>
<GID>372</GID>
<name>OUT_3</name></connection>
<connection>
<GID>349</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-31.5,45,-31.5</points>
<connection>
<GID>372</GID>
<name>OUT_4</name></connection>
<connection>
<GID>349</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-28.5,45,-28.5</points>
<connection>
<GID>372</GID>
<name>OUT_7</name></connection>
<connection>
<GID>349</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-29.5,45,-29.5</points>
<connection>
<GID>372</GID>
<name>OUT_6</name></connection>
<connection>
<GID>349</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-35.5,39,-35.5</points>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-35.5,30.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-32.5,87,-32.5</points>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection>
<connection>
<GID>367</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32,-46.5,-27.5,-46.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-44.5,-27.5,-42.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-42.5,-27.5,-42.5</points>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-28,-6,-20</points>
<connection>
<GID>347</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-28,-6,-28</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37,-29,-13,-29</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-34 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-34,-29,-34,-26.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-9,-6,-1</points>
<connection>
<GID>347</GID>
<name>load</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-34,-20.5,-34,-1</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34,-1,-6,-1</points>
<intersection>-34 1</intersection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-120,-4.5,-118</points>
<intersection>-120 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-118,12,-118</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-120,-4.5,-120</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-118,12,-95</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-118 1</intersection></vsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-117,-4.5,-94</points>
<intersection>-117 1</intersection>
<intersection>-96 2</intersection>
<intersection>-94 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-117,12,-117</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-96,-4.5,-96</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-94,12,-94</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-118,-4.5,-116</points>
<intersection>-118 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-116,12,-116</points>
<connection>
<GID>382</GID>
<name>IN_2</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-118,-4.5,-118</points>
<connection>
<GID>387</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-116,12,-93</points>
<connection>
<GID>381</GID>
<name>IN_2</name></connection>
<intersection>-116 1</intersection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-115,-4.5,-92</points>
<intersection>-115 1</intersection>
<intersection>-94 2</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-115,12,-115</points>
<connection>
<GID>382</GID>
<name>IN_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-94,-4.5,-94</points>
<connection>
<GID>386</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-92,12,-92</points>
<connection>
<GID>381</GID>
<name>IN_3</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-116,-4.5,-114</points>
<intersection>-116 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-114,12,-114</points>
<connection>
<GID>382</GID>
<name>IN_4</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-116,-4.5,-116</points>
<connection>
<GID>387</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-114,12,-91</points>
<connection>
<GID>381</GID>
<name>IN_4</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-113,-4.5,-90</points>
<intersection>-113 1</intersection>
<intersection>-92 2</intersection>
<intersection>-90 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-113,12,-113</points>
<connection>
<GID>382</GID>
<name>IN_5</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-92,-4.5,-92</points>
<connection>
<GID>386</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-4.5,-90,12,-90</points>
<connection>
<GID>381</GID>
<name>IN_5</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-114,-4.5,-112</points>
<intersection>-114 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-112,12,-112</points>
<connection>
<GID>382</GID>
<name>IN_6</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-114,-4.5,-114</points>
<connection>
<GID>387</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-112,12,-89</points>
<connection>
<GID>381</GID>
<name>IN_6</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-111,-4.5,-88</points>
<intersection>-111 1</intersection>
<intersection>-90 2</intersection>
<intersection>-88 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-111,12,-111</points>
<connection>
<GID>382</GID>
<name>IN_7</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-90,-4.5,-90</points>
<connection>
<GID>386</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-88,12,-88</points>
<connection>
<GID>381</GID>
<name>IN_7</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-110,-4.5,-87</points>
<intersection>-110 1</intersection>
<intersection>-108 2</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-110,12,-110</points>
<connection>
<GID>382</GID>
<name>IN_8</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-108,-4.5,-108</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-87,12,-87</points>
<connection>
<GID>381</GID>
<name>IN_8</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-109,-4.5,-84</points>
<intersection>-109 1</intersection>
<intersection>-86 4</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-109,12,-109</points>
<connection>
<GID>382</GID>
<name>IN_9</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-84,-4.5,-84</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-86,12,-86</points>
<connection>
<GID>381</GID>
<name>IN_9</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-108,-4.5,-85</points>
<intersection>-108 1</intersection>
<intersection>-106 2</intersection>
<intersection>-85 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-108,12,-108</points>
<connection>
<GID>382</GID>
<name>IN_10</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-106,-4.5,-106</points>
<connection>
<GID>385</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-85,12,-85</points>
<connection>
<GID>381</GID>
<name>IN_10</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-107,-4.5,-82</points>
<intersection>-107 1</intersection>
<intersection>-84 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-107,12,-107</points>
<connection>
<GID>382</GID>
<name>IN_11</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-82,-4.5,-82</points>
<connection>
<GID>384</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-84,12,-84</points>
<connection>
<GID>381</GID>
<name>IN_11</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-106,-4.5,-83</points>
<intersection>-106 1</intersection>
<intersection>-104 2</intersection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-106,12,-106</points>
<connection>
<GID>382</GID>
<name>IN_12</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-104,-4.5,-104</points>
<connection>
<GID>385</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-83,12,-83</points>
<connection>
<GID>381</GID>
<name>IN_12</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-105,-4.5,-80</points>
<intersection>-105 1</intersection>
<intersection>-82 3</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-105,12,-105</points>
<connection>
<GID>382</GID>
<name>IN_13</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-80,-4.5,-80</points>
<connection>
<GID>384</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-82,12,-82</points>
<connection>
<GID>381</GID>
<name>IN_13</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-104,-4.5,-81</points>
<intersection>-104 1</intersection>
<intersection>-102 2</intersection>
<intersection>-81 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-104,12,-104</points>
<connection>
<GID>382</GID>
<name>IN_14</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-102,-4.5,-102</points>
<connection>
<GID>385</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-81,12,-81</points>
<connection>
<GID>381</GID>
<name>IN_14</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-103,-4.5,-78</points>
<intersection>-103 1</intersection>
<intersection>-80 3</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-103,12,-103</points>
<connection>
<GID>382</GID>
<name>IN_15</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-78,-4.5,-78</points>
<connection>
<GID>384</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-80,12,-80</points>
<connection>
<GID>381</GID>
<name>IN_15</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-69.5,2.5,-69.5</points>
<connection>
<GID>392</GID>
<name>ENABLE</name></connection>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-64,54,-64</points>
<intersection>-2 8</intersection>
<intersection>54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>54,-115.5,54,-64</points>
<intersection>-115.5 18</intersection>
<intersection>-110.5 19</intersection>
<intersection>-105.5 20</intersection>
<intersection>-100.5 21</intersection>
<intersection>-95.5 22</intersection>
<intersection>-90.5 23</intersection>
<intersection>-85.5 24</intersection>
<intersection>-80.5 25</intersection>
<intersection>-64 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-2,-72.5,-2,-64</points>
<intersection>-72.5 10</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-2,-72.5,2.5,-72.5</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-2 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>54,-115.5,57,-115.5</points>
<connection>
<GID>420</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>54,-110.5,57,-110.5</points>
<connection>
<GID>419</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>54,-105.5,57,-105.5</points>
<connection>
<GID>418</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>54,-100.5,57,-100.5</points>
<connection>
<GID>417</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>54,-95.5,57,-95.5</points>
<connection>
<GID>416</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>54,-90.5,57,-90.5</points>
<connection>
<GID>415</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>54,-85.5,57,-85.5</points>
<connection>
<GID>414</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>54,-80.5,57,-80.5</points>
<connection>
<GID>413</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-101.5,9.5,-72.5</points>
<intersection>-101.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-72.5,9.5,-72.5</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-101.5,14,-101.5</points>
<connection>
<GID>382</GID>
<name>ENABLE_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-78.5,14,-71.5</points>
<connection>
<GID>381</GID>
<name>ENABLE_0</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-71.5,14,-71.5</points>
<connection>
<GID>392</GID>
<name>OUT_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-114.5,30.5,-114.5</points>
<connection>
<GID>397</GID>
<name>carry_out</name></connection>
<connection>
<GID>398</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-118,17.5,-101.5</points>
<intersection>-118 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-101.5,27.5,-101.5</points>
<connection>
<GID>397</GID>
<name>IN_B_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-118,17.5,-118</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-116,18,-102.5</points>
<intersection>-116 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-102.5,27.5,-102.5</points>
<connection>
<GID>397</GID>
<name>IN_B_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-116,18,-116</points>
<connection>
<GID>382</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-114,18.5,-103.5</points>
<intersection>-114 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-103.5,27.5,-103.5</points>
<connection>
<GID>397</GID>
<name>IN_B_2</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-114,18.5,-114</points>
<connection>
<GID>382</GID>
<name>OUT_4</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-112,19,-104.5</points>
<intersection>-112 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-104.5,27.5,-104.5</points>
<connection>
<GID>397</GID>
<name>IN_B_3</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-112,19,-112</points>
<connection>
<GID>382</GID>
<name>OUT_6</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-117.5,21,-110</points>
<intersection>-117.5 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-117.5,27.5,-117.5</points>
<connection>
<GID>398</GID>
<name>IN_B_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-110,21,-110</points>
<connection>
<GID>382</GID>
<name>OUT_8</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-118.5,20.5,-108</points>
<intersection>-118.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-118.5,27.5,-118.5</points>
<connection>
<GID>398</GID>
<name>IN_B_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-108,20.5,-108</points>
<connection>
<GID>382</GID>
<name>OUT_10</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-119.5,20,-106</points>
<intersection>-119.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-119.5,27.5,-119.5</points>
<connection>
<GID>398</GID>
<name>IN_B_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-106,20,-106</points>
<connection>
<GID>382</GID>
<name>OUT_12</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-120.5,19.5,-104</points>
<intersection>-120.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-120.5,27.5,-120.5</points>
<connection>
<GID>398</GID>
<name>IN_B_3</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-104,19.5,-104</points>
<connection>
<GID>382</GID>
<name>OUT_14</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-117,21.5,-108.5</points>
<intersection>-117 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-108.5,27.5,-108.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-117,21.5,-117</points>
<connection>
<GID>382</GID>
<name>OUT_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-115,21.5,-109.5</points>
<intersection>-115 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-109.5,27.5,-109.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-115,21.5,-115</points>
<connection>
<GID>382</GID>
<name>OUT_3</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-113,21.5,-110.5</points>
<intersection>-113 2</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-110.5,27.5,-110.5</points>
<connection>
<GID>397</GID>
<name>IN_2</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-113,21.5,-113</points>
<connection>
<GID>382</GID>
<name>OUT_5</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-111.5,21.5,-111</points>
<intersection>-111.5 1</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-111.5,27.5,-111.5</points>
<connection>
<GID>397</GID>
<name>IN_3</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-111,21.5,-111</points>
<connection>
<GID>382</GID>
<name>OUT_7</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-124.5,23.5,-109</points>
<intersection>-124.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-124.5,27.5,-124.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-109,23.5,-109</points>
<connection>
<GID>382</GID>
<name>OUT_9</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-125.5,23,-107</points>
<intersection>-125.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-125.5,27.5,-125.5</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-107,23,-107</points>
<connection>
<GID>382</GID>
<name>OUT_11</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-126.5,22.5,-105</points>
<intersection>-126.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-126.5,27.5,-126.5</points>
<connection>
<GID>398</GID>
<name>IN_2</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-105,22.5,-105</points>
<connection>
<GID>382</GID>
<name>OUT_13</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-127.5,22,-103</points>
<intersection>-127.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-127.5,27.5,-127.5</points>
<connection>
<GID>398</GID>
<name>IN_3</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-103,22,-103</points>
<connection>
<GID>382</GID>
<name>OUT_15</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-97,17,-95</points>
<intersection>-97 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-97,24,-97</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-95,17,-95</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-95,24,-95</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-95,16,-94</points>
<connection>
<GID>381</GID>
<name>OUT_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-93.5,19.5,-93</points>
<intersection>-93.5 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-93.5,29,-93.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-93,19.5,-93</points>
<connection>
<GID>381</GID>
<name>OUT_2</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-91.5,29,-91.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-92,16,-91.5</points>
<connection>
<GID>381</GID>
<name>OUT_3</name></connection>
<intersection>-91.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-90,24,-90</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-91,16,-90</points>
<connection>
<GID>381</GID>
<name>OUT_4</name></connection>
<intersection>-90 1</intersection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-90,17,-88</points>
<intersection>-90 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-88,24,-88</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-90,17,-90</points>
<connection>
<GID>381</GID>
<name>OUT_5</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-89,18,-86.5</points>
<intersection>-89 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-86.5,29,-86.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-89,18,-89</points>
<connection>
<GID>381</GID>
<name>OUT_6</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-88,17.5,-84.5</points>
<intersection>-88 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-84.5,29,-84.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-88,17.5,-88</points>
<connection>
<GID>381</GID>
<name>OUT_7</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-87,17,-83</points>
<intersection>-87 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-83,24,-83</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-87,17,-87</points>
<connection>
<GID>381</GID>
<name>OUT_8</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-86,17,-81</points>
<intersection>-86 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-81,24,-81</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-86,17,-86</points>
<connection>
<GID>381</GID>
<name>OUT_9</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-85,17.5,-79.5</points>
<intersection>-85 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-79.5,29,-79.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-85,17.5,-85</points>
<connection>
<GID>381</GID>
<name>OUT_10</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-84,17.5,-77.5</points>
<intersection>-84 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-77.5,29,-77.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-84,17.5,-84</points>
<connection>
<GID>381</GID>
<name>OUT_11</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-83,17,-76</points>
<intersection>-83 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-76,24,-76</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-83,17,-83</points>
<connection>
<GID>381</GID>
<name>OUT_12</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-82,17,-74</points>
<intersection>-82 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-74,24,-74</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-82,17,-82</points>
<connection>
<GID>381</GID>
<name>OUT_13</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-81,16.5,-72.5</points>
<intersection>-81 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-72.5,29,-72.5</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-81,16.5,-81</points>
<connection>
<GID>381</GID>
<name>OUT_14</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-80,16,-70.5</points>
<connection>
<GID>381</GID>
<name>OUT_15</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-70.5,29,-70.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-119,45,-105</points>
<intersection>-119 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-119,55,-119</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-105,45,-105</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-114,45,-106</points>
<intersection>-114 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-114,55,-114</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-106,45,-106</points>
<connection>
<GID>397</GID>
<name>OUT_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-109,45,-107</points>
<intersection>-109 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-109,55,-109</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-107,45,-107</points>
<connection>
<GID>397</GID>
<name>OUT_2</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-108,45,-104</points>
<intersection>-108 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-104,55,-104</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-108,45,-108</points>
<connection>
<GID>397</GID>
<name>OUT_3</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-121,45,-99</points>
<intersection>-121 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-99,55,-99</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-121,45,-121</points>
<connection>
<GID>398</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-122,45,-94</points>
<intersection>-122 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-94,55,-94</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-122,45,-122</points>
<connection>
<GID>398</GID>
<name>OUT_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-123,45,-89</points>
<intersection>-123 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-89,55,-89</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-123,45,-123</points>
<connection>
<GID>398</GID>
<name>OUT_2</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-124,45,-84</points>
<intersection>-124 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-84,55,-84</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-124,45,-124</points>
<connection>
<GID>398</GID>
<name>OUT_3</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-117,42.5,-96</points>
<intersection>-117 1</intersection>
<intersection>-96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-117,55,-117</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-96,42.5,-96</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-112,45,-92.5</points>
<intersection>-112 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-92.5,45,-92.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-112,55,-112</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-107,42.5,-89</points>
<intersection>-107 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-89,42.5,-89</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-107,55,-107</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-102,45,-85.5</points>
<intersection>-102 2</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-85.5,45,-85.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-102,55,-102</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-97,42.5,-82</points>
<intersection>-97 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-82,42.5,-82</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-97,55,-97</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-92,45,-78.5</points>
<intersection>-92 2</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-78.5,45,-78.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-92,55,-92</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-87,42.5,-75</points>
<intersection>-87 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-75,42.5,-75</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-87,55,-87</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-82,45,-71.5</points>
<intersection>-82 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-71.5,45,-71.5</points>
<connection>
<GID>412</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-82,55,-82</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-118,66.5,-103</points>
<intersection>-118 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-103,74.5,-103</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection>
<intersection>67.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-118,66.5,-118</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>67.5,-108.5,67.5,-103</points>
<intersection>-108.5 8</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>67.5,-108.5,88.5,-108.5</points>
<intersection>67.5 7</intersection>
<intersection>88.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>88.5,-109,88.5,-108.5</points>
<connection>
<GID>431</GID>
<name>N_in2</name></connection>
<intersection>-108.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-113,66.5,-102</points>
<intersection>-113 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-102,74.5,-102</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection>
<intersection>68 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-113,66.5,-113</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>68,-108,68,-102</points>
<intersection>-108 8</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68,-108,86,-108</points>
<intersection>68 7</intersection>
<intersection>86 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>86,-109,86,-108</points>
<connection>
<GID>430</GID>
<name>N_in2</name></connection>
<intersection>-108 8</intersection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-108,66.5,-101</points>
<intersection>-108 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-101,74.5,-101</points>
<connection>
<GID>421</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection>
<intersection>68.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-108,66.5,-108</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>68.5,-107.5,68.5,-101</points>
<intersection>-107.5 8</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-107.5,83.5,-107.5</points>
<intersection>68.5 7</intersection>
<intersection>83.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>83.5,-109,83.5,-107.5</points>
<connection>
<GID>429</GID>
<name>N_in2</name></connection>
<intersection>-107.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-103,66.5,-100</points>
<intersection>-103 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-100,74.5,-100</points>
<connection>
<GID>421</GID>
<name>IN_3</name></connection>
<intersection>66.5 0</intersection>
<intersection>69 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-103,66.5,-103</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>69,-107,69,-100</points>
<intersection>-107 9</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>69,-107,81,-107</points>
<intersection>69 8</intersection>
<intersection>81 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>81,-109,81,-107</points>
<connection>
<GID>428</GID>
<name>N_in2</name></connection>
<intersection>-107 9</intersection></vsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-99,66.5,-98</points>
<intersection>-99 1</intersection>
<intersection>-98 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-99,74.5,-99</points>
<connection>
<GID>421</GID>
<name>IN_4</name></connection>
<intersection>66.5 0</intersection>
<intersection>69.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-98,66.5,-98</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>69.5,-106.5,69.5,-99</points>
<intersection>-106.5 9</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>69.5,-106.5,78.5,-106.5</points>
<intersection>69.5 8</intersection>
<intersection>78.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>78.5,-109,78.5,-106.5</points>
<connection>
<GID>427</GID>
<name>N_in2</name></connection>
<intersection>-106.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-98,66.5,-93</points>
<intersection>-98 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-98,74.5,-98</points>
<connection>
<GID>421</GID>
<name>IN_5</name></connection>
<intersection>66.5 0</intersection>
<intersection>70 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-93,66.5,-93</points>
<connection>
<GID>415</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70,-106,70,-98</points>
<intersection>-106 8</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>70,-106,76,-106</points>
<intersection>70 7</intersection>
<intersection>76 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>76,-109,76,-106</points>
<connection>
<GID>426</GID>
<name>N_in2</name></connection>
<intersection>-106 8</intersection></vsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-97,66.5,-88</points>
<intersection>-97 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-97,74.5,-97</points>
<connection>
<GID>421</GID>
<name>IN_6</name></connection>
<intersection>66.5 0</intersection>
<intersection>70.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-88,66.5,-88</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70.5,-105.5,70.5,-97</points>
<intersection>-105.5 8</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-105.5,73.5,-105.5</points>
<intersection>70.5 7</intersection>
<intersection>73.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>73.5,-109,73.5,-105.5</points>
<connection>
<GID>425</GID>
<name>N_in2</name></connection>
<intersection>-105.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-96,66.5,-83</points>
<intersection>-96 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-83,66.5,-83</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-96,74.5,-96</points>
<connection>
<GID>421</GID>
<name>IN_7</name></connection>
<intersection>66.5 0</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-109,71,-96</points>
<connection>
<GID>424</GID>
<name>N_in2</name></connection>
<intersection>-96 2</intersection></vsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-44,172,-44</points>
<connection>
<GID>479</GID>
<name>OUT_7</name></connection>
<intersection>172 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>172,-44,172,-34</points>
<intersection>-44 1</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>172,-34,185,-34</points>
<connection>
<GID>461</GID>
<name>IN_3</name></connection>
<connection>
<GID>444</GID>
<name>IN_3</name></connection>
<intersection>172 4</intersection>
<intersection>183.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>183.5,-40,183.5,-34</points>
<intersection>-40 8</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-40,185,-40</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>183.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-45,185,-45</points>
<connection>
<GID>479</GID>
<name>OUT_6</name></connection>
<connection>
<GID>462</GID>
<name>IN_3</name></connection>
<connection>
<GID>445</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-56,171,-46</points>
<intersection>-56 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-56,185,-56</points>
<connection>
<GID>463</GID>
<name>IN_3</name></connection>
<connection>
<GID>446</GID>
<name>IN_3</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-46,171,-46</points>
<connection>
<GID>479</GID>
<name>OUT_5</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-65.5,170.5,-47</points>
<intersection>-65.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-65.5,185,-65.5</points>
<connection>
<GID>464</GID>
<name>IN_3</name></connection>
<connection>
<GID>447</GID>
<name>IN_3</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-47,170.5,-47</points>
<connection>
<GID>479</GID>
<name>OUT_4</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-76.5,170,-48</points>
<intersection>-76.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-76.5,185,-76.5</points>
<connection>
<GID>465</GID>
<name>IN_3</name></connection>
<connection>
<GID>448</GID>
<name>IN_3</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-48,170,-48</points>
<connection>
<GID>479</GID>
<name>OUT_3</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-87.5,169.5,-49</points>
<intersection>-87.5 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-87.5,185,-87.5</points>
<connection>
<GID>466</GID>
<name>IN_3</name></connection>
<connection>
<GID>449</GID>
<name>IN_3</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-49,169.5,-49</points>
<connection>
<GID>479</GID>
<name>OUT_2</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-98,169,-50</points>
<intersection>-98 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169,-98,185,-98</points>
<connection>
<GID>467</GID>
<name>IN_3</name></connection>
<connection>
<GID>450</GID>
<name>IN_3</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-50,169,-50</points>
<connection>
<GID>479</GID>
<name>OUT_1</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-109,168.5,-51</points>
<intersection>-109 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-51,168.5,-51</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-109,185,-109</points>
<connection>
<GID>468</GID>
<name>IN_3</name></connection>
<connection>
<GID>451</GID>
<name>IN_3</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-57,167.5,-36</points>
<intersection>-57 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-36,185,-36</points>
<connection>
<GID>461</GID>
<name>IN_2</name></connection>
<connection>
<GID>444</GID>
<name>IN_2</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-57,167.5,-57</points>
<connection>
<GID>480</GID>
<name>OUT_7</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-58,167,-47</points>
<intersection>-58 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-47,185,-47</points>
<connection>
<GID>462</GID>
<name>IN_2</name></connection>
<connection>
<GID>445</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-58,167,-58</points>
<connection>
<GID>480</GID>
<name>OUT_6</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-59,172.5,-59</points>
<connection>
<GID>480</GID>
<name>OUT_5</name></connection>
<intersection>172.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>172.5,-59,172.5,-58</points>
<connection>
<GID>446</GID>
<name>IN_2</name></connection>
<intersection>-59 1</intersection>
<intersection>-58 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-58,185,-58</points>
<connection>
<GID>463</GID>
<name>IN_2</name></connection>
<intersection>172.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-67.5,166.5,-60</points>
<intersection>-67.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-67.5,185,-67.5</points>
<connection>
<GID>464</GID>
<name>IN_2</name></connection>
<connection>
<GID>447</GID>
<name>IN_2</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-60,166.5,-60</points>
<connection>
<GID>480</GID>
<name>OUT_4</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-78.5,166,-61</points>
<intersection>-78.5 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-78.5,185,-78.5</points>
<connection>
<GID>465</GID>
<name>IN_2</name></connection>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-61,166,-61</points>
<connection>
<GID>480</GID>
<name>OUT_3</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-89.5,165.5,-62</points>
<intersection>-89.5 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-89.5,185,-89.5</points>
<connection>
<GID>466</GID>
<name>IN_2</name></connection>
<connection>
<GID>449</GID>
<name>IN_2</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-62,165.5,-62</points>
<connection>
<GID>480</GID>
<name>OUT_2</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-100,165,-63</points>
<intersection>-100 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-63,165,-63</points>
<connection>
<GID>480</GID>
<name>OUT_1</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-100,185,-100</points>
<connection>
<GID>467</GID>
<name>IN_2</name></connection>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-111,168,-64</points>
<intersection>-111 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-111,185,-111</points>
<connection>
<GID>468</GID>
<name>IN_2</name></connection>
<connection>
<GID>451</GID>
<name>IN_2</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-64,168,-64</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-70.5,163.5,-38</points>
<intersection>-70.5 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-38,185,-38</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-70.5,163.5,-70.5</points>
<connection>
<GID>442</GID>
<name>OUT_7</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-71.5,163,-49</points>
<intersection>-71.5 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-49,185,-49</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-71.5,163,-71.5</points>
<connection>
<GID>442</GID>
<name>OUT_6</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-72.5,162.5,-60</points>
<intersection>-72.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-60,185,-60</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-72.5,162.5,-72.5</points>
<connection>
<GID>442</GID>
<name>OUT_5</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-73.5,162,-69.5</points>
<intersection>-73.5 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-69.5,185,-69.5</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-73.5,162,-73.5</points>
<connection>
<GID>442</GID>
<name>OUT_4</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-80.5,161.5,-74.5</points>
<intersection>-80.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-80.5,185,-80.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-74.5,161.5,-74.5</points>
<connection>
<GID>442</GID>
<name>OUT_3</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-91.5,161,-75.5</points>
<intersection>-91.5 1</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-91.5,185,-91.5</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-75.5,161,-75.5</points>
<connection>
<GID>442</GID>
<name>OUT_2</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-102,160.5,-76.5</points>
<intersection>-102 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-102,185,-102</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-76.5,160.5,-76.5</points>
<connection>
<GID>442</GID>
<name>OUT_1</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-113,160,-77.5</points>
<intersection>-113 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-77.5,160,-77.5</points>
<connection>
<GID>442</GID>
<name>OUT_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-113,185,-113</points>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<connection>
<GID>451</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-83.5,159,-40</points>
<intersection>-83.5 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159,-40,172.5,-40</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-83.5,159,-83.5</points>
<connection>
<GID>443</GID>
<name>OUT_7</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-84.5,158.5,-51</points>
<intersection>-84.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,-51,185,-51</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-84.5,158.5,-84.5</points>
<connection>
<GID>443</GID>
<name>OUT_6</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-85.5,158,-62</points>
<intersection>-85.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,-62,185,-62</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-85.5,158,-85.5</points>
<connection>
<GID>443</GID>
<name>OUT_5</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-71.5,185,-71.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>154 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>154,-86.5,154,-71.5</points>
<connection>
<GID>443</GID>
<name>OUT_4</name></connection>
<intersection>-71.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-87.5,157,-82.5</points>
<intersection>-87.5 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-82.5,185,-82.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-87.5,157,-87.5</points>
<connection>
<GID>443</GID>
<name>OUT_3</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-93.5,156.5,-88.5</points>
<intersection>-93.5 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-93.5,185,-93.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-88.5,156.5,-88.5</points>
<connection>
<GID>443</GID>
<name>OUT_2</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-104,156,-89.5</points>
<intersection>-104 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-104,185,-104</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-89.5,156,-89.5</points>
<connection>
<GID>443</GID>
<name>OUT_1</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-65.5,197,-37</points>
<intersection>-65.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-37,197,-37</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-65.5,202.5,-65.5</points>
<connection>
<GID>452</GID>
<name>IN_7</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-66.5,197,-48</points>
<intersection>-66.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-48,197,-48</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-66.5,202.5,-66.5</points>
<connection>
<GID>452</GID>
<name>IN_6</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-67.5,197,-59</points>
<intersection>-67.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-59,197,-59</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-67.5,202.5,-67.5</points>
<connection>
<GID>452</GID>
<name>IN_5</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>178.5,-68.5,202.5,-68.5</points>
<connection>
<GID>452</GID>
<name>IN_4</name></connection>
<connection>
<GID>447</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-79.5,197,-69.5</points>
<intersection>-79.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-79.5,197,-79.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-69.5,202.5,-69.5</points>
<connection>
<GID>452</GID>
<name>IN_3</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-90.5,197,-70.5</points>
<intersection>-90.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-90.5,197,-90.5</points>
<connection>
<GID>449</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-70.5,202.5,-70.5</points>
<connection>
<GID>452</GID>
<name>IN_2</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-101,197,-71.5</points>
<intersection>-101 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-101,197,-101</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-71.5,202.5,-71.5</points>
<connection>
<GID>452</GID>
<name>IN_1</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-112,197,-72.5</points>
<intersection>-112 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-72.5,202.5,-72.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-112,197,-112</points>
<connection>
<GID>451</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-115,155.5,-90.5</points>
<intersection>-115 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-115,185,-115</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-90.5,155.5,-90.5</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-96,145.5,-53</points>
<intersection>-96 10</intersection>
<intersection>-92.5 8</intersection>
<intersection>-79.5 7</intersection>
<intersection>-66 6</intersection>
<intersection>-53 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>145.5,-53,149,-53</points>
<connection>
<GID>479</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>145.5,-66,149,-66</points>
<connection>
<GID>480</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>145.5,-79.5,149,-79.5</points>
<connection>
<GID>442</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>145.5,-92.5,149,-92.5</points>
<connection>
<GID>443</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>142.5,-96,145.5,-96</points>
<connection>
<GID>454</GID>
<name>CLK</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-107,176.5,-29</points>
<connection>
<GID>451</GID>
<name>SEL_0</name></connection>
<connection>
<GID>450</GID>
<name>SEL_0</name></connection>
<connection>
<GID>449</GID>
<name>SEL_0</name></connection>
<connection>
<GID>448</GID>
<name>SEL_0</name></connection>
<connection>
<GID>447</GID>
<name>SEL_0</name></connection>
<connection>
<GID>446</GID>
<name>SEL_0</name></connection>
<connection>
<GID>445</GID>
<name>SEL_0</name></connection>
<connection>
<GID>444</GID>
<name>SEL_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-29,176.5,-29</points>
<intersection>123 2</intersection>
<intersection>176.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-55,123,-29</points>
<intersection>-55 3</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-55,123,-55</points>
<connection>
<GID>453</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-107,175.5,-29.5</points>
<connection>
<GID>451</GID>
<name>SEL_1</name></connection>
<connection>
<GID>450</GID>
<name>SEL_1</name></connection>
<connection>
<GID>449</GID>
<name>SEL_1</name></connection>
<connection>
<GID>448</GID>
<name>SEL_1</name></connection>
<connection>
<GID>447</GID>
<name>SEL_1</name></connection>
<connection>
<GID>446</GID>
<name>SEL_1</name></connection>
<connection>
<GID>445</GID>
<name>SEL_1</name></connection>
<connection>
<GID>444</GID>
<name>SEL_1</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-29.5,175.5,-29.5</points>
<intersection>122.5 2</intersection>
<intersection>175.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>122.5,-53,122.5,-29.5</points>
<intersection>-53 3</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-53,122.5,-53</points>
<connection>
<GID>453</GID>
<name>OUT_1</name></connection>
<intersection>122.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-76.5,191.5,-37</points>
<intersection>-76.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-37,191.5,-37</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-76.5,202.5,-76.5</points>
<connection>
<GID>469</GID>
<name>IN_7</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-77.5,191.5,-48</points>
<intersection>-77.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-48,191.5,-48</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-77.5,202.5,-77.5</points>
<connection>
<GID>469</GID>
<name>IN_6</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-78.5,191.5,-59</points>
<intersection>-78.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-59,191.5,-59</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-78.5,202.5,-78.5</points>
<connection>
<GID>469</GID>
<name>IN_5</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-79.5,191.5,-68.5</points>
<intersection>-79.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-68.5,191.5,-68.5</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-79.5,202.5,-79.5</points>
<connection>
<GID>469</GID>
<name>IN_4</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-80.5,202.5,-80.5</points>
<connection>
<GID>469</GID>
<name>IN_3</name></connection>
<intersection>191.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>191.5,-80.5,191.5,-79.5</points>
<intersection>-80.5 1</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-79.5,191.5,-79.5</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>191.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-90.5,191.5,-81.5</points>
<intersection>-90.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-90.5,191.5,-90.5</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-81.5,202.5,-81.5</points>
<connection>
<GID>469</GID>
<name>IN_2</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-101,191.5,-82.5</points>
<intersection>-101 1</intersection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-101,191.5,-101</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-82.5,202.5,-82.5</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-112,191.5,-83.5</points>
<intersection>-112 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-83.5,202.5,-83.5</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-112,191.5,-112</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-107,189,-30.5</points>
<connection>
<GID>468</GID>
<name>SEL_0</name></connection>
<connection>
<GID>467</GID>
<name>SEL_0</name></connection>
<connection>
<GID>466</GID>
<name>SEL_0</name></connection>
<connection>
<GID>465</GID>
<name>SEL_0</name></connection>
<connection>
<GID>464</GID>
<name>SEL_0</name></connection>
<connection>
<GID>463</GID>
<name>SEL_0</name></connection>
<connection>
<GID>462</GID>
<name>SEL_0</name></connection>
<connection>
<GID>461</GID>
<name>SEL_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-30.5,189,-30.5</points>
<intersection>124 2</intersection>
<intersection>189 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-69,124,-30.5</points>
<intersection>-69 3</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-69,124,-69</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-107,188,-30</points>
<connection>
<GID>468</GID>
<name>SEL_1</name></connection>
<connection>
<GID>467</GID>
<name>SEL_1</name></connection>
<connection>
<GID>466</GID>
<name>SEL_1</name></connection>
<connection>
<GID>465</GID>
<name>SEL_1</name></connection>
<connection>
<GID>464</GID>
<name>SEL_1</name></connection>
<connection>
<GID>463</GID>
<name>SEL_1</name></connection>
<connection>
<GID>462</GID>
<name>SEL_1</name></connection>
<connection>
<GID>461</GID>
<name>SEL_1</name></connection>
<intersection>-30 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>123.5,-30,188,-30</points>
<intersection>123.5 16</intersection>
<intersection>188 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>123.5,-67,123.5,-30</points>
<intersection>-67 18</intersection>
<intersection>-30 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>122,-67,123.5,-67</points>
<connection>
<GID>460</GID>
<name>OUT_1</name></connection>
<intersection>123.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-83.5,144.5,-44</points>
<intersection>-83.5 6</intersection>
<intersection>-70.5 3</intersection>
<intersection>-62.5 4</intersection>
<intersection>-57 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-44,146,-44</points>
<connection>
<GID>479</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-57,146,-57</points>
<connection>
<GID>480</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144.5,-70.5,146,-70.5</points>
<connection>
<GID>442</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>138,-62.5,144.5,-62.5</points>
<connection>
<GID>471</GID>
<name>OUT_3</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>144.5,-83.5,146,-83.5</points>
<connection>
<GID>443</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-84.5,144,-45</points>
<intersection>-84.5 6</intersection>
<intersection>-71.5 5</intersection>
<intersection>-64.5 2</intersection>
<intersection>-58 3</intersection>
<intersection>-45 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-64.5,144,-64.5</points>
<connection>
<GID>471</GID>
<name>OUT_2</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144,-58,146,-58</points>
<connection>
<GID>480</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>144,-45,146,-45</points>
<connection>
<GID>479</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>144,-71.5,146,-71.5</points>
<connection>
<GID>442</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>144,-84.5,146,-84.5</points>
<connection>
<GID>443</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-85.5,143.5,-46</points>
<intersection>-85.5 6</intersection>
<intersection>-72.5 3</intersection>
<intersection>-66.5 2</intersection>
<intersection>-59 4</intersection>
<intersection>-46 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-66.5,143.5,-66.5</points>
<connection>
<GID>471</GID>
<name>OUT_1</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>143.5,-72.5,146,-72.5</points>
<connection>
<GID>442</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>143.5,-59,146,-59</points>
<connection>
<GID>480</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>143.5,-46,146,-46</points>
<connection>
<GID>479</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>143.5,-85.5,146,-85.5</points>
<connection>
<GID>443</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-86.5,143,-47</points>
<intersection>-86.5 6</intersection>
<intersection>-73.5 3</intersection>
<intersection>-68.5 2</intersection>
<intersection>-60 4</intersection>
<intersection>-47 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-68.5,143,-68.5</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>143,-73.5,146,-73.5</points>
<connection>
<GID>442</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>143,-60,146,-60</points>
<connection>
<GID>480</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>143,-47,146,-47</points>
<connection>
<GID>479</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>143,-86.5,146,-86.5</points>
<connection>
<GID>443</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-87.5,142.5,-48</points>
<intersection>-87.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-61 3</intersection>
<intersection>-48 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-74.5,146,-74.5</points>
<connection>
<GID>472</GID>
<name>OUT_3</name></connection>
<connection>
<GID>442</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>142.5,-61,146,-61</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142.5,-48,146,-48</points>
<connection>
<GID>479</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>142.5,-87.5,146,-87.5</points>
<connection>
<GID>443</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-88.5,142,-49</points>
<intersection>-88.5 5</intersection>
<intersection>-76.5 2</intersection>
<intersection>-75.5 4</intersection>
<intersection>-62 3</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-49,146,-49</points>
<connection>
<GID>479</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-76.5,142,-76.5</points>
<connection>
<GID>472</GID>
<name>OUT_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>142,-62,146,-62</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142,-75.5,146,-75.5</points>
<connection>
<GID>442</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>142,-88.5,146,-88.5</points>
<connection>
<GID>443</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-89.5,141.5,-50</points>
<intersection>-89.5 5</intersection>
<intersection>-78.5 2</intersection>
<intersection>-76.5 4</intersection>
<intersection>-63 3</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-50,146,-50</points>
<connection>
<GID>479</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-78.5,141.5,-78.5</points>
<connection>
<GID>472</GID>
<name>OUT_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141.5,-63,146,-63</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,-76.5,146,-76.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>141.5,-89.5,146,-89.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-90.5,141,-51</points>
<intersection>-90.5 5</intersection>
<intersection>-80.5 2</intersection>
<intersection>-77.5 4</intersection>
<intersection>-64 3</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-51,146,-51</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-80.5,141,-80.5</points>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141,-64,146,-64</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141,-77.5,146,-77.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>141,-90.5,146,-90.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-42,148,-34</points>
<intersection>-42 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-34,148,-34</points>
<connection>
<GID>474</GID>
<name>OUT_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-42,149,-42</points>
<connection>
<GID>479</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-55,148,-33</points>
<intersection>-55 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-33,148,-33</points>
<connection>
<GID>474</GID>
<name>OUT_1</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-55,149,-55</points>
<connection>
<GID>480</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-68.5,148,-32</points>
<intersection>-68.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-32,148,-32</points>
<connection>
<GID>474</GID>
<name>OUT_2</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-68.5,149,-68.5</points>
<connection>
<GID>442</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-81.5,148,-31</points>
<intersection>-81.5 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-31,148,-31</points>
<connection>
<GID>474</GID>
<name>OUT_3</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-81.5,149,-81.5</points>
<connection>
<GID>443</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-32,132,-32</points>
<connection>
<GID>475</GID>
<name>OUT_0</name></connection>
<intersection>132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132,-32,132,-31</points>
<connection>
<GID>474</GID>
<name>ENABLE</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-48,136.5,-37</points>
<intersection>-48 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-37,136.5,-37</points>
<intersection>131.5 3</intersection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-48,136.5,-48</points>
<connection>
<GID>477</GID>
<name>OUT_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-37,131.5,-34</points>
<intersection>-37 1</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>131.5,-34,132,-34</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>131.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-46,137,-36.5</points>
<intersection>-46 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-36.5,137,-36.5</points>
<intersection>132 3</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-46,137,-46</points>
<connection>
<GID>477</GID>
<name>OUT_1</name></connection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132,-36.5,132,-33</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire></page 4>
<page 5>
<PageViewport>-224.059,164.368,1553.94,-752.632</PageViewport>
<gate>
<ID>582</ID>
<type>AA_LABEL</type>
<position>50.5,-56.5</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>583</ID>
<type>AA_INVERTER</type>
<position>-1.5,-21.5</position>
<input>
<ID>IN_0</ID>751 </input>
<output>
<ID>OUT_0</ID>752 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_TOGGLE</type>
<position>23,3</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_LABEL</type>
<position>0.5,-29</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>AA_LABEL</type>
<position>0.5,-30.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>587</ID>
<type>AE_REGISTER8</type>
<position>27.5,-13</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>690 </input>
<input>
<ID>IN_2</ID>691 </input>
<input>
<ID>IN_3</ID>692 </input>
<input>
<ID>IN_4</ID>693 </input>
<input>
<ID>IN_5</ID>694 </input>
<input>
<ID>IN_6</ID>695 </input>
<input>
<ID>IN_7</ID>696 </input>
<output>
<ID>OUT_0</ID>704 </output>
<output>
<ID>OUT_1</ID>703 </output>
<output>
<ID>OUT_2</ID>702 </output>
<output>
<ID>OUT_3</ID>701 </output>
<output>
<ID>OUT_4</ID>700 </output>
<output>
<ID>OUT_5</ID>699 </output>
<output>
<ID>OUT_6</ID>698 </output>
<output>
<ID>OUT_7</ID>697 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>750 </input>
<input>
<ID>count_enable</ID>712 </input>
<input>
<ID>count_up</ID>712 </input>
<input>
<ID>load</ID>752 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_REGISTER8</type>
<position>44.5,-13</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>703 </input>
<input>
<ID>IN_2</ID>702 </input>
<input>
<ID>IN_3</ID>701 </input>
<input>
<ID>IN_4</ID>700 </input>
<input>
<ID>IN_5</ID>699 </input>
<input>
<ID>IN_6</ID>698 </input>
<input>
<ID>IN_7</ID>697 </input>
<output>
<ID>OUT_0</ID>715 </output>
<output>
<ID>OUT_1</ID>714 </output>
<output>
<ID>OUT_2</ID>710 </output>
<output>
<ID>OUT_3</ID>709 </output>
<output>
<ID>OUT_4</ID>708 </output>
<output>
<ID>OUT_5</ID>707 </output>
<output>
<ID>OUT_6</ID>706 </output>
<output>
<ID>OUT_7</ID>705 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>711 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-72.5</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>939 </output>
<output>
<ID>OUT_1</ID>938 </output>
<output>
<ID>OUT_2</ID>937 </output>
<output>
<ID>OUT_3</ID>936 </output>
<output>
<ID>OUT_4</ID>935 </output>
<output>
<ID>OUT_5</ID>934 </output>
<output>
<ID>OUT_6</ID>933 </output>
<output>
<ID>OUT_7</ID>932 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>993 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 169</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_REGISTER8</type>
<position>82.5,-51.5</position>
<input>
<ID>IN_0</ID>739 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>741 </input>
<input>
<ID>IN_3</ID>742 </input>
<input>
<ID>IN_4</ID>743 </input>
<input>
<ID>IN_5</ID>738 </input>
<input>
<ID>IN_6</ID>745 </input>
<input>
<ID>IN_7</ID>744 </input>
<output>
<ID>OUT_0</ID>723 </output>
<output>
<ID>OUT_1</ID>722 </output>
<output>
<ID>OUT_2</ID>721 </output>
<output>
<ID>OUT_3</ID>720 </output>
<output>
<ID>OUT_4</ID>719 </output>
<output>
<ID>OUT_5</ID>718 </output>
<output>
<ID>OUT_6</ID>717 </output>
<output>
<ID>OUT_7</ID>716 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>713 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-85.5</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>947 </output>
<output>
<ID>OUT_1</ID>946 </output>
<output>
<ID>OUT_2</ID>945 </output>
<output>
<ID>OUT_3</ID>944 </output>
<output>
<ID>OUT_4</ID>943 </output>
<output>
<ID>OUT_5</ID>942 </output>
<output>
<ID>OUT_6</ID>941 </output>
<output>
<ID>OUT_7</ID>940 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>994 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 147</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>590</ID>
<type>AE_RAM_8x8</type>
<position>59.5,-12.5</position>
<input>
<ID>ADDRESS_0</ID>715 </input>
<input>
<ID>ADDRESS_1</ID>714 </input>
<input>
<ID>ADDRESS_2</ID>710 </input>
<input>
<ID>ADDRESS_3</ID>709 </input>
<input>
<ID>ADDRESS_4</ID>708 </input>
<input>
<ID>ADDRESS_5</ID>707 </input>
<input>
<ID>ADDRESS_6</ID>706 </input>
<input>
<ID>ADDRESS_7</ID>705 </input>
<input>
<ID>DATA_IN_0</ID>746 </input>
<input>
<ID>DATA_IN_1</ID>731 </input>
<input>
<ID>DATA_IN_2</ID>732 </input>
<input>
<ID>DATA_IN_3</ID>733 </input>
<input>
<ID>DATA_IN_4</ID>734 </input>
<input>
<ID>DATA_IN_5</ID>735 </input>
<input>
<ID>DATA_IN_6</ID>736 </input>
<input>
<ID>DATA_IN_7</ID>737 </input>
<output>
<ID>DATA_OUT_0</ID>746 </output>
<output>
<ID>DATA_OUT_1</ID>731 </output>
<output>
<ID>DATA_OUT_2</ID>732 </output>
<output>
<ID>DATA_OUT_3</ID>733 </output>
<output>
<ID>DATA_OUT_4</ID>734 </output>
<output>
<ID>DATA_OUT_5</ID>735 </output>
<output>
<ID>DATA_OUT_6</ID>736 </output>
<output>
<ID>DATA_OUT_7</ID>737 </output>
<input>
<ID>ENABLE_0</ID>730 </input>
<input>
<ID>write_enable</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>591</ID>
<type>AE_REGISTER8</type>
<position>100,-51.5</position>
<input>
<ID>IN_0</ID>723 </input>
<input>
<ID>IN_1</ID>722 </input>
<input>
<ID>IN_2</ID>721 </input>
<input>
<ID>IN_3</ID>720 </input>
<input>
<ID>IN_4</ID>719 </input>
<input>
<ID>IN_5</ID>718 </input>
<input>
<ID>IN_6</ID>717 </input>
<input>
<ID>IN_7</ID>716 </input>
<output>
<ID>OUT_0</ID>725 </output>
<output>
<ID>OUT_1</ID>726 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>724 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>592</ID>
<type>DD_KEYPAD_HEX</type>
<position>8,-19</position>
<output>
<ID>OUT_0</ID>689 </output>
<output>
<ID>OUT_1</ID>690 </output>
<output>
<ID>OUT_2</ID>691 </output>
<output>
<ID>OUT_3</ID>692 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>593</ID>
<type>DD_KEYPAD_HEX</type>
<position>8,-7</position>
<output>
<ID>OUT_0</ID>693 </output>
<output>
<ID>OUT_1</ID>694 </output>
<output>
<ID>OUT_2</ID>695 </output>
<output>
<ID>OUT_3</ID>696 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>594</ID>
<type>BB_CLOCK</type>
<position>-3.5,-44.5</position>
<output>
<ID>CLK</ID>748 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>595</ID>
<type>AA_TOGGLE</type>
<position>25.5,6</position>
<output>
<ID>OUT_0</ID>712 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_LABEL</type>
<position>13,4</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>597</ID>
<type>AA_LABEL</type>
<position>13,6.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>598</ID>
<type>AA_TOGGLE</type>
<position>38.5,3.5</position>
<output>
<ID>OUT_0</ID>711 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_TOGGLE</type>
<position>26.5,-41.5</position>
<output>
<ID>OUT_0</ID>728 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_LABEL</type>
<position>21,-38.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>601</ID>
<type>AA_TOGGLE</type>
<position>79.5,-59.5</position>
<output>
<ID>OUT_0</ID>713 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>602</ID>
<type>AA_LABEL</type>
<position>22.5,-5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>603</ID>
<type>AA_LABEL</type>
<position>39,-5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>604</ID>
<type>AA_LABEL</type>
<position>59.5,-4</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>605</ID>
<type>AA_LABEL</type>
<position>86.5,-59</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>606</ID>
<type>AA_TOGGLE</type>
<position>96.5,-59.5</position>
<output>
<ID>OUT_0</ID>724 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>607</ID>
<type>BE_ROM_8x8</type>
<position>112.5,-51</position>
<input>
<ID>ADDRESS_0</ID>725 </input>
<input>
<ID>ADDRESS_1</ID>726 </input>
<input>
<ID>ENABLE_0</ID>747 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_TOGGLE</type>
<position>69.5,-10</position>
<output>
<ID>OUT_0</ID>729 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_TOGGLE</type>
<position>69.5,-13</position>
<output>
<ID>OUT_0</ID>730 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_LABEL</type>
<position>76,-9.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>611</ID>
<type>AA_LABEL</type>
<position>76.5,-12.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>612</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>73,-51</position>
<input>
<ID>ENABLE_0</ID>730 </input>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>731 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>733 </input>
<input>
<ID>IN_4</ID>734 </input>
<input>
<ID>IN_5</ID>735 </input>
<input>
<ID>IN_6</ID>736 </input>
<input>
<ID>IN_7</ID>737 </input>
<output>
<ID>OUT_0</ID>739 </output>
<output>
<ID>OUT_1</ID>740 </output>
<output>
<ID>OUT_2</ID>741 </output>
<output>
<ID>OUT_3</ID>742 </output>
<output>
<ID>OUT_4</ID>743 </output>
<output>
<ID>OUT_5</ID>738 </output>
<output>
<ID>OUT_6</ID>745 </output>
<output>
<ID>OUT_7</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>613</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>51,-51</position>
<input>
<ID>ENABLE_0</ID>729 </input>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>962 </input>
<input>
<ID>IN_2</ID>961 </input>
<input>
<ID>IN_3</ID>960 </input>
<input>
<ID>IN_4</ID>959 </input>
<input>
<ID>IN_5</ID>958 </input>
<input>
<ID>IN_6</ID>957 </input>
<input>
<ID>IN_7</ID>956 </input>
<output>
<ID>OUT_0</ID>746 </output>
<output>
<ID>OUT_1</ID>731 </output>
<output>
<ID>OUT_2</ID>732 </output>
<output>
<ID>OUT_3</ID>733 </output>
<output>
<ID>OUT_4</ID>734 </output>
<output>
<ID>OUT_5</ID>735 </output>
<output>
<ID>OUT_6</ID>736 </output>
<output>
<ID>OUT_7</ID>737 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>614</ID>
<type>AA_LABEL</type>
<position>101.5,-58.5</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>615</ID>
<type>AA_TOGGLE</type>
<position>121.5,-30.5</position>
<output>
<ID>OUT_0</ID>747 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_LABEL</type>
<position>123,-27.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>22.5,-26</position>
<input>
<ID>IN_0</ID>727 </input>
<input>
<ID>IN_1</ID>751 </input>
<output>
<ID>OUT</ID>750 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_AND2</type>
<position>8,-43.5</position>
<input>
<ID>IN_0</ID>749 </input>
<input>
<ID>IN_1</ID>748 </input>
<output>
<ID>OUT</ID>727 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_TOGGLE</type>
<position>2.5,-40.5</position>
<output>
<ID>OUT_0</ID>749 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>620</ID>
<type>AA_TOGGLE</type>
<position>-6.5,-27</position>
<output>
<ID>OUT_0</ID>751 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>621</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>46.5,-85.5</position>
<input>
<ID>ENABLE_0</ID>772 </input>
<input>
<ID>IN_0</ID>1004 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1010 </input>
<input>
<ID>IN_11</ID>1017 </input>
<input>
<ID>IN_12</ID>1012 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1013 </input>
<input>
<ID>IN_15</ID>1019 </input>
<input>
<ID>IN_2</ID>1006 </input>
<input>
<ID>IN_3</ID>1007 </input>
<input>
<ID>IN_4</ID>1008 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1009 </input>
<input>
<ID>IN_7</ID>1015 </input>
<input>
<ID>IN_8</ID>1010 </input>
<input>
<ID>IN_9</ID>1016 </input>
<output>
<ID>OUT_0</ID>790 </output>
<output>
<ID>OUT_1</ID>791 </output>
<output>
<ID>OUT_10</ID>800 </output>
<output>
<ID>OUT_11</ID>801 </output>
<output>
<ID>OUT_12</ID>802 </output>
<output>
<ID>OUT_13</ID>803 </output>
<output>
<ID>OUT_14</ID>804 </output>
<output>
<ID>OUT_15</ID>805 </output>
<output>
<ID>OUT_2</ID>792 </output>
<output>
<ID>OUT_3</ID>793 </output>
<output>
<ID>OUT_4</ID>794 </output>
<output>
<ID>OUT_5</ID>795 </output>
<output>
<ID>OUT_6</ID>796 </output>
<output>
<ID>OUT_7</ID>797 </output>
<output>
<ID>OUT_8</ID>798 </output>
<output>
<ID>OUT_9</ID>799 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>622</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>46.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>771 </input>
<input>
<ID>IN_0</ID>1004 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1011 </input>
<input>
<ID>IN_11</ID>1017 </input>
<input>
<ID>IN_12</ID>1012 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1013 </input>
<input>
<ID>IN_15</ID>1019 </input>
<input>
<ID>IN_2</ID>1006 </input>
<input>
<ID>IN_3</ID>1007 </input>
<input>
<ID>IN_4</ID>1008 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1009 </input>
<input>
<ID>IN_7</ID>1015 </input>
<input>
<ID>IN_8</ID>1010 </input>
<input>
<ID>IN_9</ID>1016 </input>
<output>
<ID>OUT_0</ID>774 </output>
<output>
<ID>OUT_1</ID>782 </output>
<output>
<ID>OUT_10</ID>779 </output>
<output>
<ID>OUT_11</ID>787 </output>
<output>
<ID>OUT_12</ID>780 </output>
<output>
<ID>OUT_13</ID>788 </output>
<output>
<ID>OUT_14</ID>781 </output>
<output>
<ID>OUT_15</ID>789 </output>
<output>
<ID>OUT_2</ID>775 </output>
<output>
<ID>OUT_3</ID>783 </output>
<output>
<ID>OUT_4</ID>776 </output>
<output>
<ID>OUT_5</ID>784 </output>
<output>
<ID>OUT_6</ID>777 </output>
<output>
<ID>OUT_7</ID>785 </output>
<output>
<ID>OUT_8</ID>778 </output>
<output>
<ID>OUT_9</ID>786 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_LABEL</type>
<position>24,-72.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>626</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-99</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>955 </output>
<output>
<ID>OUT_1</ID>954 </output>
<output>
<ID>OUT_2</ID>953 </output>
<output>
<ID>OUT_3</ID>952 </output>
<output>
<ID>OUT_4</ID>951 </output>
<output>
<ID>OUT_5</ID>950 </output>
<output>
<ID>OUT_6</ID>949 </output>
<output>
<ID>OUT_7</ID>948 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>995 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-112</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>971 </output>
<output>
<ID>OUT_1</ID>962 </output>
<output>
<ID>OUT_2</ID>961 </output>
<output>
<ID>OUT_3</ID>960 </output>
<output>
<ID>OUT_4</ID>959 </output>
<output>
<ID>OUT_5</ID>958 </output>
<output>
<ID>OUT_6</ID>957 </output>
<output>
<ID>OUT_7</ID>956 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>996 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_MUX_4x1</type>
<position>-50,-61.5</position>
<input>
<ID>IN_0</ID>956 </input>
<input>
<ID>IN_1</ID>948 </input>
<input>
<ID>IN_2</ID>940 </input>
<input>
<ID>IN_3</ID>932 </input>
<output>
<ID>OUT</ID>963 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>629</ID>
<type>AE_MUX_4x1</type>
<position>-50,-72.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>949 </input>
<input>
<ID>IN_2</ID>941 </input>
<input>
<ID>IN_3</ID>933 </input>
<output>
<ID>OUT</ID>964 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_MUX_4x1</type>
<position>-50,-83.5</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>950 </input>
<input>
<ID>IN_2</ID>942 </input>
<input>
<ID>IN_3</ID>934 </input>
<output>
<ID>OUT</ID>965 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>631</ID>
<type>AE_MUX_4x1</type>
<position>-50,-93</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>951 </input>
<input>
<ID>IN_2</ID>943 </input>
<input>
<ID>IN_3</ID>935 </input>
<output>
<ID>OUT</ID>966 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>632</ID>
<type>AE_MUX_4x1</type>
<position>-50,-104</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>952 </input>
<input>
<ID>IN_2</ID>944 </input>
<input>
<ID>IN_3</ID>936 </input>
<output>
<ID>OUT</ID>967 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>633</ID>
<type>AE_MUX_4x1</type>
<position>-50,-115</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>953 </input>
<input>
<ID>IN_2</ID>945 </input>
<input>
<ID>IN_3</ID>937 </input>
<output>
<ID>OUT</ID>968 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>634</ID>
<type>AE_MUX_4x1</type>
<position>-50,-125.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>954 </input>
<input>
<ID>IN_2</ID>946 </input>
<input>
<ID>IN_3</ID>938 </input>
<output>
<ID>OUT</ID>969 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>635</ID>
<type>AE_MUX_4x1</type>
<position>-50,-136.5</position>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>955 </input>
<input>
<ID>IN_2</ID>947 </input>
<input>
<ID>IN_3</ID>939 </input>
<output>
<ID>OUT</ID>970 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>636</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-11.5,-94.5</position>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>969 </input>
<input>
<ID>IN_2</ID>968 </input>
<input>
<ID>IN_3</ID>967 </input>
<input>
<ID>IN_4</ID>966 </input>
<input>
<ID>IN_5</ID>965 </input>
<input>
<ID>IN_6</ID>964 </input>
<input>
<ID>IN_7</ID>963 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 147</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>637</ID>
<type>DD_KEYPAD_HEX</type>
<position>-108.5,-76.5</position>
<output>
<ID>OUT_0</ID>973 </output>
<output>
<ID>OUT_1</ID>974 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>638</ID>
<type>BB_CLOCK</type>
<position>-87,-120.5</position>
<output>
<ID>CLK</ID>972 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_LABEL</type>
<position>-75,-105</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>640</ID>
<type>AA_LABEL</type>
<position>-75,-91.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>641</ID>
<type>AA_LABEL</type>
<position>-75,-78.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>642</ID>
<type>AA_LABEL</type>
<position>-75,-65</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>643</ID>
<type>AA_LABEL</type>
<position>-110,-69.5</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>644</ID>
<type>DD_KEYPAD_HEX</type>
<position>-108.5,-90.5</position>
<output>
<ID>OUT_0</ID>983 </output>
<output>
<ID>OUT_1</ID>984 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-61.5</position>
<input>
<ID>IN_0</ID>932 </input>
<input>
<ID>IN_1</ID>948 </input>
<input>
<ID>IN_2</ID>940 </input>
<input>
<ID>IN_3</ID>932 </input>
<output>
<ID>OUT</ID>975 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-72.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>949 </input>
<input>
<ID>IN_2</ID>941 </input>
<input>
<ID>IN_3</ID>933 </input>
<output>
<ID>OUT</ID>976 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-83.5</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>950 </input>
<input>
<ID>IN_2</ID>942 </input>
<input>
<ID>IN_3</ID>934 </input>
<output>
<ID>OUT</ID>977 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>648</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-93</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>951 </input>
<input>
<ID>IN_2</ID>943 </input>
<input>
<ID>IN_3</ID>935 </input>
<output>
<ID>OUT</ID>978 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-104</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>952 </input>
<input>
<ID>IN_2</ID>944 </input>
<input>
<ID>IN_3</ID>936 </input>
<output>
<ID>OUT</ID>979 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-115</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>953 </input>
<input>
<ID>IN_2</ID>945 </input>
<input>
<ID>IN_3</ID>937 </input>
<output>
<ID>OUT</ID>980 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>651</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-125.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>954 </input>
<input>
<ID>IN_2</ID>946 </input>
<input>
<ID>IN_3</ID>938 </input>
<output>
<ID>OUT</ID>981 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>652</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-136.5</position>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>955 </input>
<input>
<ID>IN_2</ID>947 </input>
<input>
<ID>IN_3</ID>939 </input>
<output>
<ID>OUT</ID>982 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>653</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-9.5,-105</position>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>980 </input>
<input>
<ID>IN_3</ID>979 </input>
<input>
<ID>IN_4</ID>978 </input>
<input>
<ID>IN_5</ID>977 </input>
<input>
<ID>IN_6</ID>976 </input>
<input>
<ID>IN_7</ID>975 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 169</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>654</ID>
<type>AA_LABEL</type>
<position>-110,-83.5</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>655</ID>
<type>DD_KEYPAD_HEX</type>
<position>-92.5,-90</position>
<output>
<ID>OUT_0</ID>988 </output>
<output>
<ID>OUT_1</ID>987 </output>
<output>
<ID>OUT_2</ID>986 </output>
<output>
<ID>OUT_3</ID>985 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>656</ID>
<type>DD_KEYPAD_HEX</type>
<position>-92.5,-102</position>
<output>
<ID>OUT_0</ID>992 </output>
<output>
<ID>OUT_1</ID>991 </output>
<output>
<ID>OUT_2</ID>990 </output>
<output>
<ID>OUT_3</ID>989 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_LABEL</type>
<position>-92.5,-83</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>658</ID>
<type>BA_DECODER_2x4</type>
<position>-90.5,-57</position>
<input>
<ID>ENABLE</ID>997 </input>
<input>
<ID>IN_0</ID>998 </input>
<input>
<ID>IN_1</ID>999 </input>
<output>
<ID>OUT_0</ID>993 </output>
<output>
<ID>OUT_1</ID>994 </output>
<output>
<ID>OUT_2</ID>995 </output>
<output>
<ID>OUT_3</ID>996 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_TOGGLE</type>
<position>-96.5,-56.5</position>
<output>
<ID>OUT_0</ID>997 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_LABEL</type>
<position>-99,-55</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>661</ID>
<type>DD_KEYPAD_HEX</type>
<position>-95.5,-69.5</position>
<output>
<ID>OUT_0</ID>998 </output>
<output>
<ID>OUT_1</ID>999 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_LABEL</type>
<position>-95,-62.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>668</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>6.5,-83.5</position>
<input>
<ID>ENABLE_0</ID>1000 </input>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>969 </input>
<input>
<ID>IN_2</ID>968 </input>
<input>
<ID>IN_3</ID>967 </input>
<input>
<ID>IN_4</ID>966 </input>
<input>
<ID>IN_5</ID>965 </input>
<input>
<ID>IN_6</ID>964 </input>
<input>
<ID>IN_7</ID>963 </input>
<output>
<ID>OUT_0</ID>1005 </output>
<output>
<ID>OUT_1</ID>1007 </output>
<output>
<ID>OUT_2</ID>1014 </output>
<output>
<ID>OUT_3</ID>1015 </output>
<output>
<ID>OUT_4</ID>1016 </output>
<output>
<ID>OUT_5</ID>1017 </output>
<output>
<ID>OUT_6</ID>1018 </output>
<output>
<ID>OUT_7</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>670</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>6.5,-115</position>
<input>
<ID>ENABLE_0</ID>1002 </input>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>980 </input>
<input>
<ID>IN_3</ID>979 </input>
<input>
<ID>IN_4</ID>978 </input>
<input>
<ID>IN_5</ID>977 </input>
<input>
<ID>IN_6</ID>976 </input>
<input>
<ID>IN_7</ID>975 </input>
<output>
<ID>OUT_0</ID>1004 </output>
<output>
<ID>OUT_1</ID>1006 </output>
<output>
<ID>OUT_2</ID>1008 </output>
<output>
<ID>OUT_3</ID>1009 </output>
<output>
<ID>OUT_4</ID>1010 </output>
<output>
<ID>OUT_5</ID>1011 </output>
<output>
<ID>OUT_6</ID>1012 </output>
<output>
<ID>OUT_7</ID>1013 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>672</ID>
<type>EE_VDD</type>
<position>6.5,-71.5</position>
<output>
<ID>OUT_0</ID>1000 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>482</ID>
<type>AA_LABEL</type>
<position>-18.5,-88</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>675</ID>
<type>AA_LABEL</type>
<position>4,-74.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>676</ID>
<type>AA_LABEL</type>
<position>6.5,-121</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>484</ID>
<type>AA_LABEL</type>
<position>-18.5,-99</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>678</ID>
<type>EE_VDD</type>
<position>6.5,-100</position>
<output>
<ID>OUT_0</ID>1002 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>492</ID>
<type>BA_DECODER_2x4</type>
<position>38,-69</position>
<input>
<ID>ENABLE</ID>769 </input>
<input>
<ID>IN_0</ID>770 </input>
<output>
<ID>OUT_0</ID>771 </output>
<output>
<ID>OUT_1</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_TOGGLE</type>
<position>33,-67.5</position>
<output>
<ID>OUT_0</ID>769 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_TOGGLE</type>
<position>28.5,-70.5</position>
<output>
<ID>OUT_0</ID>770 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_LABEL</type>
<position>33.5,-64.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>496</ID>
<type>AA_LABEL</type>
<position>22,-70</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>497</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64,-104.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>783 </input>
<input>
<ID>IN_2</ID>784 </input>
<input>
<ID>IN_3</ID>785 </input>
<input>
<ID>IN_B_0</ID>774 </input>
<input>
<ID>IN_B_1</ID>775 </input>
<input>
<ID>IN_B_2</ID>776 </input>
<input>
<ID>IN_B_3</ID>777 </input>
<output>
<ID>OUT_0</ID>806 </output>
<output>
<ID>OUT_1</ID>807 </output>
<output>
<ID>OUT_2</ID>808 </output>
<output>
<ID>OUT_3</ID>809 </output>
<output>
<ID>carry_out</ID>773 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64,-120.5</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>787 </input>
<input>
<ID>IN_2</ID>788 </input>
<input>
<ID>IN_3</ID>789 </input>
<input>
<ID>IN_B_0</ID>778 </input>
<input>
<ID>IN_B_1</ID>779 </input>
<input>
<ID>IN_B_2</ID>780 </input>
<input>
<ID>IN_B_3</ID>781 </input>
<output>
<ID>OUT_0</ID>810 </output>
<output>
<ID>OUT_1</ID>811 </output>
<output>
<ID>OUT_2</ID>812 </output>
<output>
<ID>OUT_3</ID>813 </output>
<input>
<ID>carry_in</ID>773 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_LABEL</type>
<position>71.5,-97</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>500</ID>
<type>AA_LABEL</type>
<position>72,-125.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>501</ID>
<type>AA_LABEL</type>
<position>57.5,-98</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>502</ID>
<type>AA_LABEL</type>
<position>58,-104.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>503</ID>
<type>AA_LABEL</type>
<position>57.5,-114</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>504</ID>
<type>AA_LABEL</type>
<position>58.5,-121</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>AA_AND2</type>
<position>59.5,-94</position>
<input>
<ID>IN_0</ID>791 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_AND2</type>
<position>64.5,-90.5</position>
<input>
<ID>IN_0</ID>793 </input>
<input>
<ID>IN_1</ID>792 </input>
<output>
<ID>OUT</ID>815 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_AND2</type>
<position>59.5,-87</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>794 </input>
<output>
<ID>OUT</ID>816 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_AND2</type>
<position>64.5,-83.5</position>
<input>
<ID>IN_0</ID>797 </input>
<input>
<ID>IN_1</ID>796 </input>
<output>
<ID>OUT</ID>817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>59.5,-80</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>798 </input>
<output>
<ID>OUT</ID>818 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_AND2</type>
<position>64.5,-76.5</position>
<input>
<ID>IN_0</ID>801 </input>
<input>
<ID>IN_1</ID>800 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_AND2</type>
<position>59.5,-73</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>802 </input>
<output>
<ID>OUT</ID>820 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>64.5,-69.5</position>
<input>
<ID>IN_0</ID>805 </input>
<input>
<ID>IN_1</ID>804 </input>
<output>
<ID>OUT</ID>821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-81</position>
<input>
<ID>IN_0</ID>813 </input>
<input>
<ID>IN_1</ID>821 </input>
<output>
<ID>OUT</ID>829 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-86</position>
<input>
<ID>IN_0</ID>812 </input>
<input>
<ID>IN_1</ID>820 </input>
<output>
<ID>OUT</ID>828 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-91</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>819 </input>
<output>
<ID>OUT</ID>827 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-96</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>818 </input>
<output>
<ID>OUT</ID>826 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>517</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-101</position>
<input>
<ID>IN_0</ID>809 </input>
<input>
<ID>IN_1</ID>817 </input>
<output>
<ID>OUT</ID>825 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-106</position>
<input>
<ID>IN_0</ID>808 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>824 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-111</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>815 </input>
<output>
<ID>OUT</ID>823 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-116</position>
<input>
<ID>IN_0</ID>806 </input>
<input>
<ID>IN_1</ID>814 </input>
<output>
<ID>OUT</ID>822 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>521</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>112,-98</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>823 </input>
<input>
<ID>IN_2</ID>824 </input>
<input>
<ID>IN_3</ID>825 </input>
<input>
<ID>IN_4</ID>826 </input>
<input>
<ID>IN_5</ID>827 </input>
<input>
<ID>IN_6</ID>828 </input>
<input>
<ID>IN_7</ID>829 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 60</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_LABEL</type>
<position>89.5,-119.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>523</ID>
<type>AA_LABEL</type>
<position>90.5,-77</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>524</ID>
<type>GA_LED</type>
<position>103.5,-108</position>
<input>
<ID>N_in2</ID>829 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>525</ID>
<type>GA_LED</type>
<position>106,-108</position>
<input>
<ID>N_in2</ID>828 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>526</ID>
<type>GA_LED</type>
<position>108.5,-108</position>
<input>
<ID>N_in2</ID>827 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>527</ID>
<type>GA_LED</type>
<position>111,-108</position>
<input>
<ID>N_in2</ID>826 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>528</ID>
<type>GA_LED</type>
<position>113.5,-108</position>
<input>
<ID>N_in2</ID>825 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>529</ID>
<type>GA_LED</type>
<position>116,-108</position>
<input>
<ID>N_in2</ID>824 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>530</ID>
<type>GA_LED</type>
<position>118.5,-108</position>
<input>
<ID>N_in2</ID>823 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>531</ID>
<type>GA_LED</type>
<position>121,-108</position>
<input>
<ID>N_in2</ID>822 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>532</ID>
<type>AA_LABEL</type>
<position>121,-110</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>533</ID>
<type>AA_LABEL</type>
<position>118.5,-110</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>534</ID>
<type>AA_LABEL</type>
<position>116,-110</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>535</ID>
<type>AA_LABEL</type>
<position>113.5,-110</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>536</ID>
<type>AA_LABEL</type>
<position>111,-110</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>537</ID>
<type>AA_LABEL</type>
<position>108.5,-110</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>AA_LABEL</type>
<position>106,-110</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>539</ID>
<type>AA_LABEL</type>
<position>103.5,-110</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-115.5,53.5,-108</points>
<intersection>-115.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-115.5,60,-115.5</points>
<connection>
<GID>498</GID>
<name>IN_B_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-108,53.5,-108</points>
<connection>
<GID>622</GID>
<name>OUT_8</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-116.5,53,-106</points>
<intersection>-116.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-116.5,60,-116.5</points>
<connection>
<GID>498</GID>
<name>IN_B_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-106,53,-106</points>
<connection>
<GID>622</GID>
<name>OUT_10</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-117.5,52.5,-104</points>
<intersection>-117.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-117.5,60,-117.5</points>
<connection>
<GID>498</GID>
<name>IN_B_2</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-104,52.5,-104</points>
<connection>
<GID>622</GID>
<name>OUT_12</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-118.5,52,-102</points>
<intersection>-118.5 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-118.5,60,-118.5</points>
<connection>
<GID>498</GID>
<name>IN_B_3</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-102,52,-102</points>
<connection>
<GID>622</GID>
<name>OUT_14</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-115,54,-106.5</points>
<intersection>-115 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-106.5,60,-106.5</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-115,54,-115</points>
<connection>
<GID>622</GID>
<name>OUT_1</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-113,54,-107.5</points>
<intersection>-113 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-107.5,60,-107.5</points>
<connection>
<GID>497</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-113,54,-113</points>
<connection>
<GID>622</GID>
<name>OUT_3</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-111,54,-108.5</points>
<intersection>-111 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-108.5,60,-108.5</points>
<connection>
<GID>497</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-111,54,-111</points>
<connection>
<GID>622</GID>
<name>OUT_5</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-109.5,54,-109</points>
<intersection>-109.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-109.5,60,-109.5</points>
<connection>
<GID>497</GID>
<name>IN_3</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-109,54,-109</points>
<connection>
<GID>622</GID>
<name>OUT_7</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-122.5,56,-107</points>
<intersection>-122.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-122.5,60,-122.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-107,56,-107</points>
<connection>
<GID>622</GID>
<name>OUT_9</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-123.5,55.5,-105</points>
<intersection>-123.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-123.5,60,-123.5</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-105,55.5,-105</points>
<connection>
<GID>622</GID>
<name>OUT_11</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-124.5,55,-103</points>
<intersection>-124.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-124.5,60,-124.5</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-103,55,-103</points>
<connection>
<GID>622</GID>
<name>OUT_13</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-125.5,54.5,-101</points>
<intersection>-125.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-125.5,60,-125.5</points>
<connection>
<GID>498</GID>
<name>IN_3</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-101,54.5,-101</points>
<connection>
<GID>622</GID>
<name>OUT_15</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-95,49.5,-93</points>
<intersection>-95 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-95,56.5,-95</points>
<connection>
<GID>505</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-93,49.5,-93</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-93,56.5,-93</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-93,48.5,-92</points>
<connection>
<GID>621</GID>
<name>OUT_1</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-91.5,52,-91</points>
<intersection>-91.5 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-91.5,61.5,-91.5</points>
<connection>
<GID>506</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-91,52,-91</points>
<connection>
<GID>621</GID>
<name>OUT_2</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-89.5,61.5,-89.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-90,48.5,-89.5</points>
<connection>
<GID>621</GID>
<name>OUT_3</name></connection>
<intersection>-89.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-88,56.5,-88</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-89,48.5,-88</points>
<connection>
<GID>621</GID>
<name>OUT_4</name></connection>
<intersection>-88 1</intersection></vsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-88,49.5,-86</points>
<intersection>-88 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-86,56.5,-86</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-88,49.5,-88</points>
<connection>
<GID>621</GID>
<name>OUT_5</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-87,50.5,-84.5</points>
<intersection>-87 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-84.5,61.5,-84.5</points>
<connection>
<GID>508</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-87,50.5,-87</points>
<connection>
<GID>621</GID>
<name>OUT_6</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-86,50,-82.5</points>
<intersection>-86 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-82.5,61.5,-82.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-86,50,-86</points>
<connection>
<GID>621</GID>
<name>OUT_7</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-85,49.5,-81</points>
<intersection>-85 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-81,56.5,-81</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-85,49.5,-85</points>
<connection>
<GID>621</GID>
<name>OUT_8</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-84,49.5,-79</points>
<intersection>-84 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-79,56.5,-79</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-84,49.5,-84</points>
<connection>
<GID>621</GID>
<name>OUT_9</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-83,50,-77.5</points>
<intersection>-83 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-77.5,61.5,-77.5</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-83,50,-83</points>
<connection>
<GID>621</GID>
<name>OUT_10</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-82,50,-75.5</points>
<intersection>-82 2</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-75.5,61.5,-75.5</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-82,50,-82</points>
<connection>
<GID>621</GID>
<name>OUT_11</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-81,49.5,-74</points>
<intersection>-81 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-74,56.5,-74</points>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-81,49.5,-81</points>
<connection>
<GID>621</GID>
<name>OUT_12</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-80,49.5,-72</points>
<intersection>-80 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-72,56.5,-72</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-80,49.5,-80</points>
<connection>
<GID>621</GID>
<name>OUT_13</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-79,49,-70.5</points>
<intersection>-79 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-70.5,61.5,-70.5</points>
<connection>
<GID>512</GID>
<name>IN_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-79,49,-79</points>
<connection>
<GID>621</GID>
<name>OUT_14</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-78,48.5,-68.5</points>
<connection>
<GID>621</GID>
<name>OUT_15</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-68.5,61.5,-68.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-117,77.5,-103</points>
<intersection>-117 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-117,87.5,-117</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-103,77.5,-103</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-112,77.5,-104</points>
<intersection>-112 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-112,87.5,-112</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-104,77.5,-104</points>
<connection>
<GID>497</GID>
<name>OUT_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-107,77.5,-105</points>
<intersection>-107 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-107,87.5,-107</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-105,77.5,-105</points>
<connection>
<GID>497</GID>
<name>OUT_2</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-106,77.5,-102</points>
<intersection>-106 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-102,87.5,-102</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-106,77.5,-106</points>
<connection>
<GID>497</GID>
<name>OUT_3</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-119,77.5,-97</points>
<intersection>-119 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-97,87.5,-97</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-119,77.5,-119</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-120,77.5,-92</points>
<intersection>-120 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-92,87.5,-92</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-120,77.5,-120</points>
<connection>
<GID>498</GID>
<name>OUT_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-121,77.5,-87</points>
<intersection>-121 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-87,87.5,-87</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-121,77.5,-121</points>
<connection>
<GID>498</GID>
<name>OUT_2</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-122,77.5,-82</points>
<intersection>-122 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-82,87.5,-82</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-122,77.5,-122</points>
<connection>
<GID>498</GID>
<name>OUT_3</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-115,75,-94</points>
<intersection>-115 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-115,87.5,-115</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-94,75,-94</points>
<connection>
<GID>505</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-110,77.5,-90.5</points>
<intersection>-110 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-90.5,77.5,-90.5</points>
<connection>
<GID>506</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-110,87.5,-110</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-105,75,-87</points>
<intersection>-105 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-87,75,-87</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-105,87.5,-105</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-100,77.5,-83.5</points>
<intersection>-100 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-83.5,77.5,-83.5</points>
<connection>
<GID>508</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-100,87.5,-100</points>
<connection>
<GID>517</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-95,75,-80</points>
<intersection>-95 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-80,75,-80</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-95,87.5,-95</points>
<connection>
<GID>516</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-90,77.5,-76.5</points>
<intersection>-90 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-76.5,77.5,-76.5</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-90,87.5,-90</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-85,75,-73</points>
<intersection>-85 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-73,75,-73</points>
<connection>
<GID>511</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-85,87.5,-85</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-80,77.5,-69.5</points>
<intersection>-80 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-69.5,77.5,-69.5</points>
<connection>
<GID>512</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-80,87.5,-80</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-116,99,-101</points>
<intersection>-116 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-101,107,-101</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection>
<intersection>100 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-116,99,-116</points>
<connection>
<GID>520</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>100,-106.5,100,-101</points>
<intersection>-106.5 8</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100,-106.5,121,-106.5</points>
<intersection>100 7</intersection>
<intersection>121 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>121,-107,121,-106.5</points>
<connection>
<GID>531</GID>
<name>N_in2</name></connection>
<intersection>-106.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-111,99,-100</points>
<intersection>-111 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-100,107,-100</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection>
<intersection>100.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-111,99,-111</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>100.5,-106,100.5,-100</points>
<intersection>-106 8</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100.5,-106,118.5,-106</points>
<intersection>100.5 7</intersection>
<intersection>118.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>118.5,-107,118.5,-106</points>
<connection>
<GID>530</GID>
<name>N_in2</name></connection>
<intersection>-106 8</intersection></vsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-106,99,-99</points>
<intersection>-106 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-99,107,-99</points>
<connection>
<GID>521</GID>
<name>IN_2</name></connection>
<intersection>99 0</intersection>
<intersection>101 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-106,99,-106</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>101,-105.5,101,-99</points>
<intersection>-105.5 8</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>101,-105.5,116,-105.5</points>
<intersection>101 7</intersection>
<intersection>116 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>116,-107,116,-105.5</points>
<connection>
<GID>529</GID>
<name>N_in2</name></connection>
<intersection>-105.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-101,99,-98</points>
<intersection>-101 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-98,107,-98</points>
<connection>
<GID>521</GID>
<name>IN_3</name></connection>
<intersection>99 0</intersection>
<intersection>101.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-101,99,-101</points>
<connection>
<GID>517</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>101.5,-105,101.5,-98</points>
<intersection>-105 9</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>101.5,-105,113.5,-105</points>
<intersection>101.5 8</intersection>
<intersection>113.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>113.5,-107,113.5,-105</points>
<connection>
<GID>528</GID>
<name>N_in2</name></connection>
<intersection>-105 9</intersection></vsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-97,99,-96</points>
<intersection>-97 1</intersection>
<intersection>-96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-97,107,-97</points>
<connection>
<GID>521</GID>
<name>IN_4</name></connection>
<intersection>99 0</intersection>
<intersection>102 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-96,99,-96</points>
<connection>
<GID>516</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>102,-104.5,102,-97</points>
<intersection>-104.5 9</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>102,-104.5,111,-104.5</points>
<intersection>102 8</intersection>
<intersection>111 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>111,-107,111,-104.5</points>
<connection>
<GID>527</GID>
<name>N_in2</name></connection>
<intersection>-104.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-96,99,-91</points>
<intersection>-96 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-96,107,-96</points>
<connection>
<GID>521</GID>
<name>IN_5</name></connection>
<intersection>99 0</intersection>
<intersection>102.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-91,99,-91</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>102.5,-104,102.5,-96</points>
<intersection>-104 8</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>102.5,-104,108.5,-104</points>
<intersection>102.5 7</intersection>
<intersection>108.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>108.5,-107,108.5,-104</points>
<connection>
<GID>526</GID>
<name>N_in2</name></connection>
<intersection>-104 8</intersection></vsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-95,99,-86</points>
<intersection>-95 1</intersection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-95,107,-95</points>
<connection>
<GID>521</GID>
<name>IN_6</name></connection>
<intersection>99 0</intersection>
<intersection>103 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-86,99,-86</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>103,-103.5,103,-95</points>
<intersection>-103.5 8</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>103,-103.5,106,-103.5</points>
<intersection>103 7</intersection>
<intersection>106 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>106,-107,106,-103.5</points>
<connection>
<GID>525</GID>
<name>N_in2</name></connection>
<intersection>-103.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-94,99,-81</points>
<intersection>-94 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-81,99,-81</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-94,107,-94</points>
<connection>
<GID>521</GID>
<name>IN_7</name></connection>
<intersection>99 0</intersection>
<intersection>103.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>103.5,-107,103.5,-94</points>
<connection>
<GID>524</GID>
<name>N_in2</name></connection>
<intersection>-94 2</intersection></vsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-68.5,-53.5,-68.5</points>
<connection>
<GID>202</GID>
<name>OUT_7</name></connection>
<intersection>-53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53.5,-68.5,-53.5,-58.5</points>
<intersection>-68.5 1</intersection>
<intersection>-58.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-53.5,-58.5,-40.5,-58.5</points>
<connection>
<GID>628</GID>
<name>IN_3</name></connection>
<connection>
<GID>645</GID>
<name>IN_3</name></connection>
<intersection>-53.5 4</intersection>
<intersection>-42 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-42,-64.5,-42,-58.5</points>
<intersection>-64.5 8</intersection>
<intersection>-58.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-42,-64.5,-40.5,-64.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>-42 6</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-69.5,-40.5,-69.5</points>
<connection>
<GID>202</GID>
<name>OUT_6</name></connection>
<connection>
<GID>629</GID>
<name>IN_3</name></connection>
<connection>
<GID>646</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-80.5,-54.5,-70.5</points>
<intersection>-80.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,-80.5,-40.5,-80.5</points>
<connection>
<GID>630</GID>
<name>IN_3</name></connection>
<connection>
<GID>647</GID>
<name>IN_3</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-70.5,-54.5,-70.5</points>
<connection>
<GID>202</GID>
<name>OUT_5</name></connection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-90,-55,-71.5</points>
<intersection>-90 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-90,-40.5,-90</points>
<connection>
<GID>631</GID>
<name>IN_3</name></connection>
<connection>
<GID>648</GID>
<name>IN_3</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-71.5,-55,-71.5</points>
<connection>
<GID>202</GID>
<name>OUT_4</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-101,-55.5,-72.5</points>
<intersection>-101 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-101,-40.5,-101</points>
<connection>
<GID>632</GID>
<name>IN_3</name></connection>
<connection>
<GID>649</GID>
<name>IN_3</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-72.5,-55.5,-72.5</points>
<connection>
<GID>202</GID>
<name>OUT_3</name></connection>
<intersection>-55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-112,-56,-73.5</points>
<intersection>-112 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-112,-40.5,-112</points>
<connection>
<GID>633</GID>
<name>IN_3</name></connection>
<connection>
<GID>650</GID>
<name>IN_3</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-73.5,-56,-73.5</points>
<connection>
<GID>202</GID>
<name>OUT_2</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-122.5,-56.5,-74.5</points>
<intersection>-122.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,-122.5,-40.5,-122.5</points>
<connection>
<GID>634</GID>
<name>IN_3</name></connection>
<connection>
<GID>651</GID>
<name>IN_3</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-74.5,-56.5,-74.5</points>
<connection>
<GID>202</GID>
<name>OUT_1</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-133.5,-57,-75.5</points>
<intersection>-133.5 2</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-75.5,-57,-75.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-133.5,-40.5,-133.5</points>
<connection>
<GID>635</GID>
<name>IN_3</name></connection>
<connection>
<GID>652</GID>
<name>IN_3</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-81.5,-58,-60.5</points>
<intersection>-81.5 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-60.5,-40.5,-60.5</points>
<connection>
<GID>628</GID>
<name>IN_2</name></connection>
<connection>
<GID>645</GID>
<name>IN_2</name></connection>
<intersection>-58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-81.5,-58,-81.5</points>
<connection>
<GID>203</GID>
<name>OUT_7</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-82.5,-58.5,-71.5</points>
<intersection>-82.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-71.5,-40.5,-71.5</points>
<connection>
<GID>629</GID>
<name>IN_2</name></connection>
<connection>
<GID>646</GID>
<name>IN_2</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-82.5,-58.5,-82.5</points>
<connection>
<GID>203</GID>
<name>OUT_6</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-83.5,-53,-83.5</points>
<connection>
<GID>203</GID>
<name>OUT_5</name></connection>
<intersection>-53 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-53,-83.5,-53,-82.5</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>-83.5 1</intersection>
<intersection>-82.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-53,-82.5,-40.5,-82.5</points>
<connection>
<GID>647</GID>
<name>IN_2</name></connection>
<intersection>-53 3</intersection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-92,-59,-84.5</points>
<intersection>-92 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,-92,-40.5,-92</points>
<connection>
<GID>631</GID>
<name>IN_2</name></connection>
<connection>
<GID>648</GID>
<name>IN_2</name></connection>
<intersection>-59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-84.5,-59,-84.5</points>
<connection>
<GID>203</GID>
<name>OUT_4</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-103,-59.5,-85.5</points>
<intersection>-103 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-103,-40.5,-103</points>
<connection>
<GID>632</GID>
<name>IN_2</name></connection>
<connection>
<GID>649</GID>
<name>IN_2</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-85.5,-59.5,-85.5</points>
<connection>
<GID>203</GID>
<name>OUT_3</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-114,-60,-86.5</points>
<intersection>-114 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-114,-40.5,-114</points>
<connection>
<GID>633</GID>
<name>IN_2</name></connection>
<connection>
<GID>650</GID>
<name>IN_2</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-86.5,-60,-86.5</points>
<connection>
<GID>203</GID>
<name>OUT_2</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-124.5,-60.5,-87.5</points>
<intersection>-124.5 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-87.5,-60.5,-87.5</points>
<connection>
<GID>203</GID>
<name>OUT_1</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60.5,-124.5,-40.5,-124.5</points>
<connection>
<GID>634</GID>
<name>IN_2</name></connection>
<connection>
<GID>651</GID>
<name>IN_2</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-135.5,-57.5,-88.5</points>
<intersection>-135.5 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,-135.5,-40.5,-135.5</points>
<connection>
<GID>635</GID>
<name>IN_2</name></connection>
<connection>
<GID>652</GID>
<name>IN_2</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-88.5,-57.5,-88.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-95,-62,-62.5</points>
<intersection>-95 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-62.5,-40.5,-62.5</points>
<connection>
<GID>628</GID>
<name>IN_1</name></connection>
<connection>
<GID>645</GID>
<name>IN_1</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-95,-62,-95</points>
<connection>
<GID>626</GID>
<name>OUT_7</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-96,-62.5,-73.5</points>
<intersection>-96 2</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-73.5,-40.5,-73.5</points>
<connection>
<GID>629</GID>
<name>IN_1</name></connection>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-96,-62.5,-96</points>
<connection>
<GID>626</GID>
<name>OUT_6</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-97,-63,-84.5</points>
<intersection>-97 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-84.5,-40.5,-84.5</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<connection>
<GID>647</GID>
<name>IN_1</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-97,-63,-97</points>
<connection>
<GID>626</GID>
<name>OUT_5</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-98,-63.5,-94</points>
<intersection>-98 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-94,-40.5,-94</points>
<connection>
<GID>631</GID>
<name>IN_1</name></connection>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-98,-63.5,-98</points>
<connection>
<GID>626</GID>
<name>OUT_4</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,-105,-64,-99</points>
<intersection>-105 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-105,-40.5,-105</points>
<connection>
<GID>632</GID>
<name>IN_1</name></connection>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-99,-64,-99</points>
<connection>
<GID>626</GID>
<name>OUT_3</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-116,-64.5,-100</points>
<intersection>-116 1</intersection>
<intersection>-100 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-116,-40.5,-116</points>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<connection>
<GID>650</GID>
<name>IN_1</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-100,-64.5,-100</points>
<connection>
<GID>626</GID>
<name>OUT_2</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-126.5,-65,-101</points>
<intersection>-126.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-126.5,-40.5,-126.5</points>
<connection>
<GID>634</GID>
<name>IN_1</name></connection>
<connection>
<GID>651</GID>
<name>IN_1</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-101,-65,-101</points>
<connection>
<GID>626</GID>
<name>OUT_1</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-137.5,-65.5,-102</points>
<intersection>-137.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-102,-65.5,-102</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,-137.5,-40.5,-137.5</points>
<connection>
<GID>635</GID>
<name>IN_1</name></connection>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-153,-66.5,-108</points>
<intersection>-153 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-153,-4.5,-153</points>
<intersection>-66.5 0</intersection>
<intersection>-53 5</intersection>
<intersection>-4.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-108,-66.5,-108</points>
<connection>
<GID>627</GID>
<name>OUT_7</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-4.5,-153,-4.5,-47.5</points>
<intersection>-153 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-53,-153,-53,-64.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-4.5,-47.5,49,-47.5</points>
<connection>
<GID>613</GID>
<name>IN_7</name></connection>
<intersection>-4.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-154.5,-67,-109</points>
<intersection>-154.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,-154.5,-3,-154.5</points>
<intersection>-67 0</intersection>
<intersection>-53 7</intersection>
<intersection>-40.5 8</intersection>
<intersection>-3 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-109,-67,-109</points>
<connection>
<GID>627</GID>
<name>OUT_6</name></connection>
<intersection>-67 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-3,-154.5,-3,-48.5</points>
<intersection>-154.5 1</intersection>
<intersection>-48.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-3,-48.5,49,-48.5</points>
<connection>
<GID>613</GID>
<name>IN_6</name></connection>
<intersection>-3 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-53,-154.5,-53,-75.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-40.5,-154.5,-40.5,-75.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-155.5,-67.5,-110</points>
<intersection>-155.5 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-155.5,-1.5,-155.5</points>
<intersection>-67.5 0</intersection>
<intersection>-53 8</intersection>
<intersection>-40.5 9</intersection>
<intersection>-1.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-110,-67.5,-110</points>
<connection>
<GID>627</GID>
<name>OUT_5</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1.5,-155.5,-1.5,-49.5</points>
<intersection>-155.5 1</intersection>
<intersection>-49.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1.5,-49.5,49,-49.5</points>
<connection>
<GID>613</GID>
<name>IN_5</name></connection>
<intersection>-1.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-53,-155.5,-53,-86.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>-155.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-40.5,-155.5,-40.5,-86.5</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-155.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-157.5,0,-157.5</points>
<intersection>-68 6</intersection>
<intersection>-53 13</intersection>
<intersection>-40.5 14</intersection>
<intersection>0 11</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-68,-157.5,-68,-111</points>
<intersection>-157.5 1</intersection>
<intersection>-111 15</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>0,-157.5,0,-50.5</points>
<intersection>-157.5 1</intersection>
<intersection>-50.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>0,-50.5,49,-50.5</points>
<connection>
<GID>613</GID>
<name>IN_4</name></connection>
<intersection>0 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-53,-157.5,-53,-96</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-40.5,-157.5,-40.5,-96</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-71.5,-111,-68,-111</points>
<connection>
<GID>627</GID>
<name>OUT_4</name></connection>
<intersection>-68 6</intersection></hsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-159,-68.5,-112</points>
<intersection>-159 1</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,-159,1,-159</points>
<intersection>-68.5 0</intersection>
<intersection>-53 9</intersection>
<intersection>-40.5 10</intersection>
<intersection>1 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-112,-68.5,-112</points>
<connection>
<GID>627</GID>
<name>OUT_3</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>1,-159,1,-51.5</points>
<intersection>-159 1</intersection>
<intersection>-51.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>1,-51.5,49,-51.5</points>
<connection>
<GID>613</GID>
<name>IN_3</name></connection>
<intersection>1 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-53,-159,-53,-107</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-40.5,-159,-40.5,-107</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection></vsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-160.5,-69,-113</points>
<intersection>-160.5 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-160.5,2,-160.5</points>
<intersection>-69 0</intersection>
<intersection>-53 4</intersection>
<intersection>-40.5 5</intersection>
<intersection>2 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-113,-69,-113</points>
<connection>
<GID>627</GID>
<name>OUT_2</name></connection>
<intersection>-69 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2,-160.5,2,-52.5</points>
<intersection>-160.5 1</intersection>
<intersection>-52.5 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-53,-160.5,-53,-118</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-40.5,-160.5,-40.5,-118</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>2,-52.5,49,-52.5</points>
<connection>
<GID>613</GID>
<name>IN_2</name></connection>
<intersection>2 3</intersection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-161.5,-69.5,-114</points>
<intersection>-161.5 1</intersection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-161.5,3,-161.5</points>
<intersection>-69.5 0</intersection>
<intersection>-53 8</intersection>
<intersection>-40.5 9</intersection>
<intersection>3 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-114,-69.5,-114</points>
<connection>
<GID>627</GID>
<name>OUT_1</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>3,-161.5,3,-53.5</points>
<intersection>-161.5 1</intersection>
<intersection>-53.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>3,-53.5,49,-53.5</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<intersection>3 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-53,-161.5,-53,-128.5</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>-161.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-40.5,-161.5,-40.5,-128.5</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-161.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-90.5,-28.5,-61.5</points>
<intersection>-90.5 2</intersection>
<intersection>-80 3</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-61.5,-28.5,-61.5</points>
<connection>
<GID>628</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-90.5,-16.5,-90.5</points>
<connection>
<GID>636</GID>
<name>IN_7</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,-80,4.5,-80</points>
<connection>
<GID>668</GID>
<name>IN_7</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-91.5,-28.5,-72.5</points>
<intersection>-91.5 2</intersection>
<intersection>-81 4</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-72.5,-28.5,-72.5</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-91.5,-16.5,-91.5</points>
<connection>
<GID>636</GID>
<name>IN_6</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-28.5,-81,4.5,-81</points>
<connection>
<GID>668</GID>
<name>IN_6</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-92.5,-28.5,-82</points>
<intersection>-92.5 2</intersection>
<intersection>-83.5 1</intersection>
<intersection>-82 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-83.5,-28.5,-83.5</points>
<connection>
<GID>630</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-92.5,-16.5,-92.5</points>
<connection>
<GID>636</GID>
<name>IN_5</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,-82,4.5,-82</points>
<connection>
<GID>668</GID>
<name>IN_5</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-93.5,-16.5,-93.5</points>
<connection>
<GID>636</GID>
<name>IN_4</name></connection>
<intersection>-47 6</intersection>
<intersection>-27.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-27.5,-93.5,-27.5,-83</points>
<intersection>-93.5 1</intersection>
<intersection>-83 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-27.5,-83,4.5,-83</points>
<connection>
<GID>668</GID>
<name>IN_4</name></connection>
<intersection>-27.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-47,-93.5,-47,-93</points>
<connection>
<GID>631</GID>
<name>OUT</name></connection>
<intersection>-93.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-104,-28.5,-94.5</points>
<intersection>-104 1</intersection>
<intersection>-94.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-104,-28.5,-104</points>
<connection>
<GID>632</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-94.5,-16.5,-94.5</points>
<connection>
<GID>636</GID>
<name>IN_3</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-26.5,-94.5,-26.5,-84</points>
<intersection>-94.5 2</intersection>
<intersection>-84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-26.5,-84,4.5,-84</points>
<connection>
<GID>668</GID>
<name>IN_3</name></connection>
<intersection>-26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-115,-28.5,-95.5</points>
<intersection>-115 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-115,-28.5,-115</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-95.5,-16.5,-95.5</points>
<connection>
<GID>636</GID>
<name>IN_2</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25.5,-95.5,-25.5,-85</points>
<intersection>-95.5 2</intersection>
<intersection>-85 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25.5,-85,4.5,-85</points>
<connection>
<GID>668</GID>
<name>IN_2</name></connection>
<intersection>-25.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-125.5,-28.5,-96.5</points>
<intersection>-125.5 1</intersection>
<intersection>-96.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-125.5,-28.5,-125.5</points>
<connection>
<GID>634</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-96.5,-16.5,-96.5</points>
<connection>
<GID>636</GID>
<name>IN_1</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24.5,-96.5,-24.5,-86</points>
<intersection>-96.5 2</intersection>
<intersection>-86 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-24.5,-86,4.5,-86</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<intersection>-24.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-136.5,-28.5,-97.5</points>
<intersection>-136.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28.5,-97.5,-16.5,-97.5</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-23.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-136.5,-28.5,-136.5</points>
<connection>
<GID>635</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-23.5,-97.5,-23.5,-87</points>
<intersection>-97.5 1</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-23.5,-87,4.5,-87</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-23.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,-163,-70,-115</points>
<intersection>-163 1</intersection>
<intersection>-115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70,-163,4,-163</points>
<intersection>-70 0</intersection>
<intersection>-53 14</intersection>
<intersection>-40.5 15</intersection>
<intersection>4 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-115,-70,-115</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<intersection>-70 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>4,-163,4,-54.5</points>
<intersection>-163 1</intersection>
<intersection>-54.5 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-53,-163,-53,-139.5</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>-163 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-40.5,-163,-40.5,-139.5</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>-163 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>4,-54.5,49,-54.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>4 13</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-120.5,-80,-77.5</points>
<intersection>-120.5 10</intersection>
<intersection>-117 8</intersection>
<intersection>-104 7</intersection>
<intersection>-90.5 6</intersection>
<intersection>-77.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-80,-77.5,-76.5,-77.5</points>
<connection>
<GID>202</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-80,-90.5,-76.5,-90.5</points>
<connection>
<GID>203</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-80,-104,-76.5,-104</points>
<connection>
<GID>626</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-80,-117,-76.5,-117</points>
<connection>
<GID>627</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-83,-120.5,-80,-120.5</points>
<connection>
<GID>638</GID>
<name>CLK</name></connection>
<intersection>-80 0</intersection></hsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-131.5,-49,-53.5</points>
<connection>
<GID>635</GID>
<name>SEL_0</name></connection>
<connection>
<GID>634</GID>
<name>SEL_0</name></connection>
<connection>
<GID>633</GID>
<name>SEL_0</name></connection>
<connection>
<GID>632</GID>
<name>SEL_0</name></connection>
<connection>
<GID>631</GID>
<name>SEL_0</name></connection>
<connection>
<GID>630</GID>
<name>SEL_0</name></connection>
<connection>
<GID>629</GID>
<name>SEL_0</name></connection>
<connection>
<GID>628</GID>
<name>SEL_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-102.5,-53.5,-49,-53.5</points>
<intersection>-102.5 2</intersection>
<intersection>-49 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-102.5,-79.5,-102.5,-53.5</points>
<intersection>-79.5 3</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-79.5,-102.5,-79.5</points>
<connection>
<GID>637</GID>
<name>OUT_0</name></connection>
<intersection>-102.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-131.5,-50,-54</points>
<connection>
<GID>635</GID>
<name>SEL_1</name></connection>
<connection>
<GID>634</GID>
<name>SEL_1</name></connection>
<connection>
<GID>633</GID>
<name>SEL_1</name></connection>
<connection>
<GID>632</GID>
<name>SEL_1</name></connection>
<connection>
<GID>631</GID>
<name>SEL_1</name></connection>
<connection>
<GID>630</GID>
<name>SEL_1</name></connection>
<connection>
<GID>629</GID>
<name>SEL_1</name></connection>
<connection>
<GID>628</GID>
<name>SEL_1</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,-54,-50,-54</points>
<intersection>-103 2</intersection>
<intersection>-50 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-103,-77.5,-103,-54</points>
<intersection>-77.5 3</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-77.5,-103,-77.5</points>
<connection>
<GID>637</GID>
<name>OUT_1</name></connection>
<intersection>-103 2</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-101,-34,-61.5</points>
<intersection>-101 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-61.5,-34,-61.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-101,-14.5,-101</points>
<connection>
<GID>653</GID>
<name>IN_7</name></connection>
<intersection>-34 0</intersection>
<intersection>-28 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-28,-111.5,-28,-101</points>
<intersection>-111.5 4</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-28,-111.5,4.5,-111.5</points>
<connection>
<GID>670</GID>
<name>IN_7</name></connection>
<intersection>-28 3</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-102,-34,-72.5</points>
<intersection>-102 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-72.5,-34,-72.5</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-102,-14.5,-102</points>
<connection>
<GID>653</GID>
<name>IN_6</name></connection>
<intersection>-34 0</intersection>
<intersection>-27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-112.5,-27.5,-102</points>
<intersection>-112.5 4</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-27.5,-112.5,4.5,-112.5</points>
<connection>
<GID>670</GID>
<name>IN_6</name></connection>
<intersection>-27.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-103,-34,-83.5</points>
<intersection>-103 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-83.5,-34,-83.5</points>
<connection>
<GID>647</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-103,-14.5,-103</points>
<connection>
<GID>653</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection>
<intersection>-25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25.5,-113.5,-25.5,-103</points>
<intersection>-113.5 4</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25.5,-113.5,4.5,-113.5</points>
<connection>
<GID>670</GID>
<name>IN_5</name></connection>
<intersection>-25.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-104,-34,-93</points>
<intersection>-104 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-93,-34,-93</points>
<connection>
<GID>648</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-104,-14.5,-104</points>
<connection>
<GID>653</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection>
<intersection>-24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24,-114.5,-24,-104</points>
<intersection>-114.5 4</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-24,-114.5,4.5,-114.5</points>
<connection>
<GID>670</GID>
<name>IN_4</name></connection>
<intersection>-24 3</intersection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34,-105,-14.5,-105</points>
<connection>
<GID>653</GID>
<name>IN_3</name></connection>
<intersection>-34 2</intersection>
<intersection>-22 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34,-105,-34,-104</points>
<intersection>-105 1</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-34.5,-104,-34,-104</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>-34 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22,-115.5,-22,-105</points>
<intersection>-115.5 5</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-22,-115.5,4.5,-115.5</points>
<connection>
<GID>670</GID>
<name>IN_3</name></connection>
<intersection>-22 4</intersection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-115,-34,-106</points>
<intersection>-115 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-115,-34,-115</points>
<connection>
<GID>650</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-106,-14.5,-106</points>
<connection>
<GID>653</GID>
<name>IN_2</name></connection>
<intersection>-34 0</intersection>
<intersection>-20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-20,-116.5,-20,-106</points>
<intersection>-116.5 4</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20,-116.5,4.5,-116.5</points>
<connection>
<GID>670</GID>
<name>IN_2</name></connection>
<intersection>-20 3</intersection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-125.5,-34,-107</points>
<intersection>-125.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-125.5,-34,-125.5</points>
<connection>
<GID>651</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-107,-14.5,-107</points>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<intersection>-34 0</intersection>
<intersection>-19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19,-117.5,-19,-107</points>
<intersection>-117.5 4</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-19,-117.5,4.5,-117.5</points>
<connection>
<GID>670</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-136.5,-34,-108</points>
<intersection>-136.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-108,-14.5,-108</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection>
<intersection>-18 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-136.5,-34,-136.5</points>
<connection>
<GID>652</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,-118.5,-18,-108</points>
<intersection>-118.5 4</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-18,-118.5,4.5,-118.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-131.5,-36.5,-55</points>
<connection>
<GID>652</GID>
<name>SEL_0</name></connection>
<connection>
<GID>651</GID>
<name>SEL_0</name></connection>
<connection>
<GID>650</GID>
<name>SEL_0</name></connection>
<connection>
<GID>649</GID>
<name>SEL_0</name></connection>
<connection>
<GID>648</GID>
<name>SEL_0</name></connection>
<connection>
<GID>647</GID>
<name>SEL_0</name></connection>
<connection>
<GID>646</GID>
<name>SEL_0</name></connection>
<connection>
<GID>645</GID>
<name>SEL_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-101.5,-55,-36.5,-55</points>
<intersection>-101.5 2</intersection>
<intersection>-36.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-101.5,-93.5,-101.5,-55</points>
<intersection>-93.5 3</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-93.5,-101.5,-93.5</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-131.5,-37.5,-54.5</points>
<connection>
<GID>652</GID>
<name>SEL_1</name></connection>
<connection>
<GID>651</GID>
<name>SEL_1</name></connection>
<connection>
<GID>650</GID>
<name>SEL_1</name></connection>
<connection>
<GID>649</GID>
<name>SEL_1</name></connection>
<connection>
<GID>648</GID>
<name>SEL_1</name></connection>
<connection>
<GID>647</GID>
<name>SEL_1</name></connection>
<connection>
<GID>646</GID>
<name>SEL_1</name></connection>
<connection>
<GID>645</GID>
<name>SEL_1</name></connection>
<intersection>-54.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-102,-54.5,-37.5,-54.5</points>
<intersection>-102 16</intersection>
<intersection>-37.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-102,-91.5,-102,-54.5</points>
<intersection>-91.5 18</intersection>
<intersection>-54.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-103.5,-91.5,-102,-91.5</points>
<connection>
<GID>644</GID>
<name>OUT_1</name></connection>
<intersection>-102 16</intersection></hsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-108,-81,-68.5</points>
<intersection>-108 6</intersection>
<intersection>-95 3</intersection>
<intersection>-87 4</intersection>
<intersection>-81.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81,-68.5,-79.5,-68.5</points>
<connection>
<GID>202</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-81,-81.5,-79.5,-81.5</points>
<connection>
<GID>203</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-81,-95,-79.5,-95</points>
<connection>
<GID>626</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-87.5,-87,-81,-87</points>
<connection>
<GID>655</GID>
<name>OUT_3</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-81,-108,-79.5,-108</points>
<connection>
<GID>627</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,-109,-81.5,-69.5</points>
<intersection>-109 6</intersection>
<intersection>-96 5</intersection>
<intersection>-89 2</intersection>
<intersection>-82.5 3</intersection>
<intersection>-69.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-89,-81.5,-89</points>
<connection>
<GID>655</GID>
<name>OUT_2</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-81.5,-82.5,-79.5,-82.5</points>
<connection>
<GID>203</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-81.5,-69.5,-79.5,-69.5</points>
<connection>
<GID>202</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-81.5,-96,-79.5,-96</points>
<connection>
<GID>626</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-81.5,-109,-79.5,-109</points>
<connection>
<GID>627</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,-110,-82,-70.5</points>
<intersection>-110 6</intersection>
<intersection>-97 3</intersection>
<intersection>-91 2</intersection>
<intersection>-83.5 4</intersection>
<intersection>-70.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-91,-82,-91</points>
<connection>
<GID>655</GID>
<name>OUT_1</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-82,-97,-79.5,-97</points>
<connection>
<GID>626</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-82,-83.5,-79.5,-83.5</points>
<connection>
<GID>203</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-82,-70.5,-79.5,-70.5</points>
<connection>
<GID>202</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-82,-110,-79.5,-110</points>
<connection>
<GID>627</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82.5,-111,-82.5,-71.5</points>
<intersection>-111 6</intersection>
<intersection>-98 3</intersection>
<intersection>-93 2</intersection>
<intersection>-84.5 4</intersection>
<intersection>-71.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-93,-82.5,-93</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-82.5,-98,-79.5,-98</points>
<connection>
<GID>626</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-82.5,-84.5,-79.5,-84.5</points>
<connection>
<GID>203</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-82.5,-71.5,-79.5,-71.5</points>
<connection>
<GID>202</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-82.5,-111,-79.5,-111</points>
<connection>
<GID>627</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,-112,-83,-72.5</points>
<intersection>-112 5</intersection>
<intersection>-99 2</intersection>
<intersection>-85.5 3</intersection>
<intersection>-72.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-99,-79.5,-99</points>
<connection>
<GID>626</GID>
<name>IN_3</name></connection>
<connection>
<GID>656</GID>
<name>OUT_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-83,-85.5,-79.5,-85.5</points>
<connection>
<GID>203</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-83,-72.5,-79.5,-72.5</points>
<connection>
<GID>202</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-83,-112,-79.5,-112</points>
<connection>
<GID>627</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83.5,-113,-83.5,-73.5</points>
<intersection>-113 5</intersection>
<intersection>-101 2</intersection>
<intersection>-100 4</intersection>
<intersection>-86.5 3</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83.5,-73.5,-79.5,-73.5</points>
<connection>
<GID>202</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-101,-83.5,-101</points>
<connection>
<GID>656</GID>
<name>OUT_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-83.5,-86.5,-79.5,-86.5</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-83.5,-100,-79.5,-100</points>
<connection>
<GID>626</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-83.5,-113,-79.5,-113</points>
<connection>
<GID>627</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-114,-84,-74.5</points>
<intersection>-114 5</intersection>
<intersection>-103 2</intersection>
<intersection>-101 4</intersection>
<intersection>-87.5 3</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84,-74.5,-79.5,-74.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-103,-84,-103</points>
<connection>
<GID>656</GID>
<name>OUT_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84,-87.5,-79.5,-87.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-101,-79.5,-101</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-84,-114,-79.5,-114</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-115,-84.5,-75.5</points>
<intersection>-115 5</intersection>
<intersection>-105 2</intersection>
<intersection>-102 4</intersection>
<intersection>-88.5 3</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,-75.5,-79.5,-75.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-105,-84.5,-105</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84.5,-88.5,-79.5,-88.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84.5,-102,-79.5,-102</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-84.5,-115,-79.5,-115</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-66.5,-77.5,-58.5</points>
<intersection>-66.5 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-58.5,-77.5,-58.5</points>
<connection>
<GID>658</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-66.5,-76.5,-66.5</points>
<connection>
<GID>202</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-79.5,-77.5,-57.5</points>
<intersection>-79.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-57.5,-77.5,-57.5</points>
<connection>
<GID>658</GID>
<name>OUT_1</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-79.5,-76.5,-79.5</points>
<connection>
<GID>203</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-93,-77.5,-56.5</points>
<intersection>-93 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-56.5,-77.5,-56.5</points>
<connection>
<GID>658</GID>
<name>OUT_2</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-93,-76.5,-93</points>
<connection>
<GID>626</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-106,-77.5,-55.5</points>
<intersection>-106 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-55.5,-77.5,-55.5</points>
<connection>
<GID>658</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-106,-76.5,-106</points>
<connection>
<GID>627</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94.5,-56.5,-93.5,-56.5</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>-93.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-93.5,-56.5,-93.5,-55.5</points>
<connection>
<GID>658</GID>
<name>ENABLE</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89,-72.5,-89,-61.5</points>
<intersection>-72.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94,-61.5,-89,-61.5</points>
<intersection>-94 3</intersection>
<intersection>-89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,-72.5,-89,-72.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>-89 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-94,-61.5,-94,-58.5</points>
<intersection>-61.5 1</intersection>
<intersection>-58.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-94,-58.5,-93.5,-58.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-94 3</intersection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,-70.5,-88.5,-61</points>
<intersection>-70.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-61,-88.5,-61</points>
<intersection>-93.5 3</intersection>
<intersection>-88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,-70.5,-88.5,-70.5</points>
<connection>
<GID>661</GID>
<name>OUT_1</name></connection>
<intersection>-88.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-93.5,-61,-93.5,-57.5</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-78.5,6.5,-72.5</points>
<connection>
<GID>668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-110,6.5,-101</points>
<connection>
<GID>670</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>678</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-118.5,30.5,-93</points>
<intersection>-118.5 1</intersection>
<intersection>-93 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-118.5,44.5,-118.5</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-93,44.5,-93</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-118.5,44.5,-116</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-118.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-115,30.5,-87</points>
<intersection>-115 1</intersection>
<intersection>-92 3</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-115,44.5,-115</points>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-87,30.5,-87</points>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-92,44.5,-92</points>
<connection>
<GID>621</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-117.5,30.5,-91</points>
<intersection>-117.5 2</intersection>
<intersection>-114 1</intersection>
<intersection>-91 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-114,44.5,-114</points>
<connection>
<GID>622</GID>
<name>IN_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-117.5,30.5,-117.5</points>
<connection>
<GID>670</GID>
<name>OUT_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-91,44.5,-91</points>
<connection>
<GID>621</GID>
<name>IN_2</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-113,30.5,-86</points>
<intersection>-113 1</intersection>
<intersection>-90 3</intersection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-113,44.5,-113</points>
<connection>
<GID>622</GID>
<name>IN_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-86,30.5,-86</points>
<connection>
<GID>668</GID>
<name>OUT_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-90,44.5,-90</points>
<connection>
<GID>621</GID>
<name>IN_3</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-116.5,30.5,-112</points>
<intersection>-116.5 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-112,44.5,-112</points>
<connection>
<GID>622</GID>
<name>IN_4</name></connection>
<intersection>30.5 0</intersection>
<intersection>39.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-116.5,30.5,-116.5</points>
<connection>
<GID>670</GID>
<name>OUT_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-112,39.5,-89</points>
<intersection>-112 1</intersection>
<intersection>-89 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39.5,-89,44.5,-89</points>
<connection>
<GID>621</GID>
<name>IN_4</name></connection>
<intersection>39.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-115.5,30.5,-110</points>
<intersection>-115.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-110,44.5,-110</points>
<connection>
<GID>622</GID>
<name>IN_6</name></connection>
<intersection>30.5 0</intersection>
<intersection>44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-115.5,30.5,-115.5</points>
<connection>
<GID>670</GID>
<name>OUT_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-110,44,-87</points>
<intersection>-110 1</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>44,-87,44.5,-87</points>
<connection>
<GID>621</GID>
<name>IN_6</name></connection>
<intersection>44 3</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-114.5,30.5,-108</points>
<intersection>-114.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-108,44.5,-108</points>
<connection>
<GID>622</GID>
<name>IN_8</name></connection>
<intersection>30.5 0</intersection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-114.5,30.5,-114.5</points>
<connection>
<GID>670</GID>
<name>OUT_4</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-108,42.5,-83</points>
<intersection>-108 1</intersection>
<intersection>-85 6</intersection>
<intersection>-83 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-83,44.5,-83</points>
<connection>
<GID>621</GID>
<name>IN_10</name></connection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>42.5,-85,44.5,-85</points>
<connection>
<GID>621</GID>
<name>IN_8</name></connection>
<intersection>42.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-113.5,30.5,-106</points>
<intersection>-113.5 2</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-106,44.5,-106</points>
<connection>
<GID>622</GID>
<name>IN_10</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-113.5,30.5,-113.5</points>
<connection>
<GID>670</GID>
<name>OUT_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-112.5,30.5,-104</points>
<intersection>-112.5 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-104,44.5,-104</points>
<connection>
<GID>622</GID>
<name>IN_12</name></connection>
<intersection>30.5 0</intersection>
<intersection>43.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-112.5,30.5,-112.5</points>
<connection>
<GID>670</GID>
<name>OUT_6</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-104,43.5,-81</points>
<intersection>-104 1</intersection>
<intersection>-81 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-81,44.5,-81</points>
<connection>
<GID>621</GID>
<name>IN_12</name></connection>
<intersection>43.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-111.5,30.5,-102</points>
<intersection>-111.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-102,44.5,-102</points>
<connection>
<GID>622</GID>
<name>IN_14</name></connection>
<intersection>30.5 0</intersection>
<intersection>38 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-111.5,30.5,-111.5</points>
<connection>
<GID>670</GID>
<name>OUT_7</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-102,38,-79</points>
<intersection>-102 1</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,-79,44.5,-79</points>
<connection>
<GID>621</GID>
<name>IN_14</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-111,30.5,-85</points>
<intersection>-111 1</intersection>
<intersection>-88 3</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-111,44.5,-111</points>
<connection>
<GID>622</GID>
<name>IN_5</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-85,30.5,-85</points>
<connection>
<GID>668</GID>
<name>OUT_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-88,44.5,-88</points>
<connection>
<GID>621</GID>
<name>IN_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-109,30.5,-84</points>
<intersection>-109 1</intersection>
<intersection>-86 3</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-109,44.5,-109</points>
<connection>
<GID>622</GID>
<name>IN_7</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-84,30.5,-84</points>
<connection>
<GID>668</GID>
<name>OUT_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-86,44.5,-86</points>
<connection>
<GID>621</GID>
<name>IN_7</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-107,30.5,-83</points>
<intersection>-107 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-107,44.5,-107</points>
<connection>
<GID>622</GID>
<name>IN_9</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-83,44.5,-83</points>
<connection>
<GID>668</GID>
<name>OUT_4</name></connection>
<intersection>30.5 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-84,44.5,-83</points>
<connection>
<GID>621</GID>
<name>IN_9</name></connection>
<intersection>-83 2</intersection></vsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-105,30.5,-82</points>
<intersection>-105 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-105,44.5,-105</points>
<connection>
<GID>622</GID>
<name>IN_11</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-82,44.5,-82</points>
<connection>
<GID>621</GID>
<name>IN_11</name></connection>
<connection>
<GID>668</GID>
<name>OUT_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-103,30.5,-80</points>
<intersection>-103 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-103,44.5,-103</points>
<connection>
<GID>622</GID>
<name>IN_13</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-80,44.5,-80</points>
<connection>
<GID>621</GID>
<name>IN_13</name></connection>
<intersection>17 4</intersection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17,-81,17,-80</points>
<intersection>-81 5</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>8.5,-81,17,-81</points>
<connection>
<GID>668</GID>
<name>OUT_6</name></connection>
<intersection>17 4</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-101,30.5,-78</points>
<intersection>-101 1</intersection>
<intersection>-79 2</intersection>
<intersection>-78 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-101,44.5,-101</points>
<connection>
<GID>622</GID>
<name>IN_15</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-79,30.5,-79</points>
<intersection>8.5 4</intersection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-78,44.5,-78</points>
<connection>
<GID>621</GID>
<name>IN_15</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-80,8.5,-79</points>
<connection>
<GID>668</GID>
<name>OUT_7</name></connection>
<intersection>-79 2</intersection></vsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-22,18,-16</points>
<intersection>-22 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-16,23.5,-16</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-22,18,-22</points>
<connection>
<GID>592</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-20,18,-15</points>
<intersection>-20 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-15,23.5,-15</points>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-20,18,-20</points>
<connection>
<GID>592</GID>
<name>OUT_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-18,18,-14</points>
<intersection>-18 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-14,23.5,-14</points>
<connection>
<GID>587</GID>
<name>IN_2</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-18,18,-18</points>
<connection>
<GID>592</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-16,18,-13</points>
<intersection>-16 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-13,23.5,-13</points>
<connection>
<GID>587</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-16,18,-16</points>
<connection>
<GID>592</GID>
<name>OUT_3</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-12,18,-10</points>
<intersection>-12 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-12,23.5,-12</points>
<connection>
<GID>587</GID>
<name>IN_4</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-10,18,-10</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-11,18,-8</points>
<intersection>-11 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-11,23.5,-11</points>
<connection>
<GID>587</GID>
<name>IN_5</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-8,18,-8</points>
<connection>
<GID>593</GID>
<name>OUT_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-10,18,-6</points>
<intersection>-10 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-10,23.5,-10</points>
<connection>
<GID>587</GID>
<name>IN_6</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-6,18,-6</points>
<connection>
<GID>593</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-9,23.5,-9</points>
<connection>
<GID>587</GID>
<name>IN_7</name></connection>
<intersection>13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-9,13,-4</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-9,40.5,-9</points>
<connection>
<GID>587</GID>
<name>OUT_7</name></connection>
<connection>
<GID>588</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-10,40.5,-10</points>
<connection>
<GID>587</GID>
<name>OUT_6</name></connection>
<connection>
<GID>588</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-11,40.5,-11</points>
<connection>
<GID>587</GID>
<name>OUT_5</name></connection>
<connection>
<GID>588</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-12,40.5,-12</points>
<connection>
<GID>587</GID>
<name>OUT_4</name></connection>
<connection>
<GID>588</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-13,40.5,-13</points>
<connection>
<GID>587</GID>
<name>OUT_3</name></connection>
<connection>
<GID>588</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-14,40.5,-14</points>
<connection>
<GID>587</GID>
<name>OUT_2</name></connection>
<connection>
<GID>588</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-15,40.5,-15</points>
<connection>
<GID>587</GID>
<name>OUT_1</name></connection>
<connection>
<GID>588</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-16,40.5,-16</points>
<connection>
<GID>587</GID>
<name>OUT_0</name></connection>
<connection>
<GID>588</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-9,54.5,-9</points>
<connection>
<GID>588</GID>
<name>OUT_7</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-10,54.5,-10</points>
<connection>
<GID>588</GID>
<name>OUT_6</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-11,54.5,-11</points>
<connection>
<GID>588</GID>
<name>OUT_5</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-12,54.5,-12</points>
<connection>
<GID>588</GID>
<name>OUT_4</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-13,54.5,-13</points>
<connection>
<GID>588</GID>
<name>OUT_3</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-14,54.5,-14</points>
<connection>
<GID>588</GID>
<name>OUT_2</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-7,43.5,3.5</points>
<connection>
<GID>588</GID>
<name>load</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,3.5,43.5,3.5</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-7,27.5,6</points>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection>
<connection>
<GID>587</GID>
<name>count_enable</name></connection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-6,28.5,-6</points>
<intersection>27.5 0</intersection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-7,28.5,-6</points>
<connection>
<GID>587</GID>
<name>count_up</name></connection>
<intersection>-6 2</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>81.5,-59.5,81.5,-45.5</points>
<connection>
<GID>601</GID>
<name>OUT_0</name></connection>
<connection>
<GID>589</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-15,54.5,-15</points>
<connection>
<GID>588</GID>
<name>OUT_1</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-16,54.5,-16</points>
<connection>
<GID>588</GID>
<name>OUT_0</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-47.5,96,-47.5</points>
<connection>
<GID>589</GID>
<name>OUT_7</name></connection>
<connection>
<GID>591</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-48.5,96,-48.5</points>
<connection>
<GID>589</GID>
<name>OUT_6</name></connection>
<connection>
<GID>591</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-49.5,96,-49.5</points>
<connection>
<GID>589</GID>
<name>OUT_5</name></connection>
<connection>
<GID>591</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-50.5,96,-50.5</points>
<connection>
<GID>589</GID>
<name>OUT_4</name></connection>
<connection>
<GID>591</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-51.5,96,-51.5</points>
<connection>
<GID>589</GID>
<name>OUT_3</name></connection>
<connection>
<GID>591</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-52.5,96,-52.5</points>
<connection>
<GID>589</GID>
<name>OUT_2</name></connection>
<connection>
<GID>591</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-53.5,96,-53.5</points>
<connection>
<GID>589</GID>
<name>OUT_1</name></connection>
<connection>
<GID>591</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-54.5,96,-54.5</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-59.5,99,-45.5</points>
<connection>
<GID>591</GID>
<name>load</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-59.5,99,-59.5</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-54.5,107.5,-54.5</points>
<connection>
<GID>591</GID>
<name>OUT_0</name></connection>
<connection>
<GID>607</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-53.5,107.5,-53.5</points>
<connection>
<GID>591</GID>
<name>OUT_1</name></connection>
<connection>
<GID>607</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-43.5,43.5,-18</points>
<connection>
<GID>588</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-43.5,99,-43.5</points>
<connection>
<GID>618</GID>
<name>OUT</name></connection>
<intersection>13.5 6</intersection>
<intersection>43.5 0</intersection>
<intersection>81.5 5</intersection>
<intersection>99 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>99,-56.5,99,-43.5</points>
<connection>
<GID>591</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>81.5,-56.5,81.5,-43.5</points>
<connection>
<GID>589</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>13.5,-43.5,13.5,-25</points>
<intersection>-43.5 1</intersection>
<intersection>-25 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13.5,-25,19.5,-25</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>13.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-41.5,28.5,-18</points>
<connection>
<GID>599</GID>
<name>OUT_0</name></connection>
<connection>
<GID>587</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-41.5,101,-41.5</points>
<intersection>28.5 0</intersection>
<intersection>45.5 3</intersection>
<intersection>83.5 7</intersection>
<intersection>101 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-41.5,45.5,-18</points>
<connection>
<GID>588</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>101,-56.5,101,-41.5</points>
<connection>
<GID>591</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>83.5,-56.5,83.5,-41.5</points>
<connection>
<GID>589</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-10,67.5,-10</points>
<connection>
<GID>608</GID>
<name>OUT_0</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-25,65.5,-10</points>
<intersection>-25 4</intersection>
<intersection>-12 7</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-25,65.5,-25</points>
<intersection>51 8</intersection>
<intersection>65.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>64.5,-12,65.5,-12</points>
<connection>
<GID>590</GID>
<name>write_enable</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>51,-46,51,-25</points>
<connection>
<GID>613</GID>
<name>ENABLE_0</name></connection>
<intersection>-25 4</intersection></vsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-13,67.5,-13</points>
<connection>
<GID>590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>609</GID>
<name>OUT_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>67.5,-25,67.5,-13</points>
<intersection>-25 6</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>67.5,-25,73,-25</points>
<intersection>67.5 5</intersection>
<intersection>73 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>73,-46,73,-25</points>
<connection>
<GID>612</GID>
<name>ENABLE_0</name></connection>
<intersection>-25 6</intersection></vsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-53.5,71,-53.5</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<connection>
<GID>613</GID>
<name>OUT_1</name></connection>
<intersection>62 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>62,-53.5,62,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-52.5,71,-52.5</points>
<connection>
<GID>612</GID>
<name>IN_2</name></connection>
<connection>
<GID>613</GID>
<name>OUT_2</name></connection>
<intersection>61 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>61,-52.5,61,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_2</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-51.5,71,-51.5</points>
<connection>
<GID>612</GID>
<name>IN_3</name></connection>
<connection>
<GID>613</GID>
<name>OUT_3</name></connection>
<intersection>60 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>60,-51.5,60,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_3</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-50.5,71,-50.5</points>
<connection>
<GID>612</GID>
<name>IN_4</name></connection>
<connection>
<GID>613</GID>
<name>OUT_4</name></connection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-50.5,59,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_4</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-49.5,71,-49.5</points>
<connection>
<GID>612</GID>
<name>IN_5</name></connection>
<connection>
<GID>613</GID>
<name>OUT_5</name></connection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-49.5,58,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_5</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-48.5,71,-48.5</points>
<connection>
<GID>612</GID>
<name>IN_6</name></connection>
<connection>
<GID>613</GID>
<name>OUT_6</name></connection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-48.5,57,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_6</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-47.5,71,-47.5</points>
<connection>
<GID>612</GID>
<name>IN_7</name></connection>
<connection>
<GID>613</GID>
<name>OUT_7</name></connection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-47.5,56,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_7</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-49.5,78.5,-49.5</points>
<connection>
<GID>589</GID>
<name>IN_5</name></connection>
<connection>
<GID>612</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-54.5,78.5,-54.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-53.5,78.5,-53.5</points>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<connection>
<GID>612</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-52.5,78.5,-52.5</points>
<connection>
<GID>589</GID>
<name>IN_2</name></connection>
<connection>
<GID>612</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-51.5,78.5,-51.5</points>
<connection>
<GID>589</GID>
<name>IN_3</name></connection>
<connection>
<GID>612</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-50.5,78.5,-50.5</points>
<connection>
<GID>589</GID>
<name>IN_4</name></connection>
<connection>
<GID>612</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-47.5,78.5,-47.5</points>
<connection>
<GID>589</GID>
<name>IN_7</name></connection>
<connection>
<GID>612</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-48.5,78.5,-48.5</points>
<connection>
<GID>589</GID>
<name>IN_6</name></connection>
<connection>
<GID>612</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-54.5,71,-54.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-54.5,63,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_0</name></connection>
<intersection>-54.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117.5,-51.5,119.5,-51.5</points>
<connection>
<GID>607</GID>
<name>ENABLE_0</name></connection>
<intersection>119.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119.5,-51.5,119.5,-30.5</points>
<connection>
<GID>615</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-44.5,5,-44.5</points>
<connection>
<GID>594</GID>
<name>CLK</name></connection>
<connection>
<GID>618</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-42.5,5,-40.5</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-40.5,5,-40.5</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-26,26.5,-18</points>
<connection>
<GID>587</GID>
<name>clock</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-26,26.5,-26</points>
<connection>
<GID>617</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,-27,19.5,-27</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>-1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-27,-1.5,-24.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-7,26.5,1</points>
<connection>
<GID>587</GID>
<name>load</name></connection>
<intersection>1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1.5,-18.5,-1.5,1</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,1,26.5,1</points>
<intersection>-1.5 1</intersection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-67.5,35,-67.5</points>
<connection>
<GID>492</GID>
<name>ENABLE</name></connection>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-62,86.5,-62</points>
<intersection>30.5 8</intersection>
<intersection>86.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>86.5,-113.5,86.5,-62</points>
<intersection>-113.5 18</intersection>
<intersection>-108.5 19</intersection>
<intersection>-103.5 20</intersection>
<intersection>-98.5 21</intersection>
<intersection>-93.5 22</intersection>
<intersection>-88.5 23</intersection>
<intersection>-83.5 24</intersection>
<intersection>-78.5 25</intersection>
<intersection>-62 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>30.5,-70.5,30.5,-62</points>
<intersection>-70.5 10</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>30.5,-70.5,35,-70.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>30.5 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>86.5,-113.5,89.5,-113.5</points>
<connection>
<GID>520</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>86.5,-108.5,89.5,-108.5</points>
<connection>
<GID>519</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>86.5,-103.5,89.5,-103.5</points>
<connection>
<GID>518</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>86.5,-98.5,89.5,-98.5</points>
<connection>
<GID>517</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>86.5,-93.5,89.5,-93.5</points>
<connection>
<GID>516</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>86.5,-88.5,89.5,-88.5</points>
<connection>
<GID>515</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>86.5,-83.5,89.5,-83.5</points>
<connection>
<GID>514</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>86.5,-78.5,89.5,-78.5</points>
<connection>
<GID>513</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-99.5,42,-70.5</points>
<intersection>-99.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-70.5,42,-70.5</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-99.5,46.5,-99.5</points>
<connection>
<GID>622</GID>
<name>ENABLE_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-76.5,46.5,-69.5</points>
<connection>
<GID>621</GID>
<name>ENABLE_0</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-69.5,46.5,-69.5</points>
<connection>
<GID>492</GID>
<name>OUT_1</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-112.5,63,-112.5</points>
<connection>
<GID>497</GID>
<name>carry_out</name></connection>
<connection>
<GID>498</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-116,50,-99.5</points>
<intersection>-116 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-99.5,60,-99.5</points>
<connection>
<GID>497</GID>
<name>IN_B_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-116,50,-116</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-114,50.5,-100.5</points>
<intersection>-114 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-100.5,60,-100.5</points>
<connection>
<GID>497</GID>
<name>IN_B_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-114,50.5,-114</points>
<connection>
<GID>622</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-112,51,-101.5</points>
<intersection>-112 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-101.5,60,-101.5</points>
<connection>
<GID>497</GID>
<name>IN_B_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-112,51,-112</points>
<connection>
<GID>622</GID>
<name>OUT_4</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-110,51.5,-102.5</points>
<intersection>-110 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-102.5,60,-102.5</points>
<connection>
<GID>497</GID>
<name>IN_B_3</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-110,51.5,-110</points>
<connection>
<GID>622</GID>
<name>OUT_6</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>486.001,-80.957,734.124,-208.926</PageViewport>
<gate>
<ID>772</ID>
<type>AA_TOGGLE</type>
<position>603,-87</position>
<output>
<ID>OUT_0</ID>1085 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>773</ID>
<type>AA_LABEL</type>
<position>624.5,-81</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>774</ID>
<type>AA_LABEL</type>
<position>596.5,-86.5</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>775</ID>
<type>AE_FULLADDER_4BIT</type>
<position>655,-121</position>
<input>
<ID>IN_0</ID>1097 </input>
<input>
<ID>IN_1</ID>1098 </input>
<input>
<ID>IN_2</ID>1099 </input>
<input>
<ID>IN_3</ID>1100 </input>
<input>
<ID>IN_B_0</ID>1089 </input>
<input>
<ID>IN_B_1</ID>1090 </input>
<input>
<ID>IN_B_2</ID>1091 </input>
<input>
<ID>IN_B_3</ID>1092 </input>
<output>
<ID>OUT_0</ID>1121 </output>
<output>
<ID>OUT_1</ID>1122 </output>
<output>
<ID>OUT_2</ID>1123 </output>
<output>
<ID>OUT_3</ID>1124 </output>
<output>
<ID>carry_out</ID>1088 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>776</ID>
<type>AE_FULLADDER_4BIT</type>
<position>655,-137</position>
<input>
<ID>IN_0</ID>1101 </input>
<input>
<ID>IN_1</ID>1102 </input>
<input>
<ID>IN_2</ID>1103 </input>
<input>
<ID>IN_3</ID>1104 </input>
<input>
<ID>IN_B_0</ID>1093 </input>
<input>
<ID>IN_B_1</ID>1094 </input>
<input>
<ID>IN_B_2</ID>1095 </input>
<input>
<ID>IN_B_3</ID>1096 </input>
<output>
<ID>OUT_0</ID>1125 </output>
<output>
<ID>OUT_1</ID>1126 </output>
<output>
<ID>OUT_2</ID>1127 </output>
<output>
<ID>OUT_3</ID>1128 </output>
<input>
<ID>carry_in</ID>1088 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_LABEL</type>
<position>662.5,-113.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>778</ID>
<type>AA_LABEL</type>
<position>663,-142</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>779</ID>
<type>AA_LABEL</type>
<position>648.5,-114.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>780</ID>
<type>AA_LABEL</type>
<position>649,-121</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>781</ID>
<type>AA_LABEL</type>
<position>648.5,-130.5</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>782</ID>
<type>AA_LABEL</type>
<position>649.5,-137.5</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>650.5,-110.5</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1105 </input>
<output>
<ID>OUT</ID>1129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AA_AND2</type>
<position>655.5,-107</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1107 </input>
<output>
<ID>OUT</ID>1130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>785</ID>
<type>AA_AND2</type>
<position>650.5,-103.5</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1109 </input>
<output>
<ID>OUT</ID>1131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>AA_AND2</type>
<position>655.5,-100</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1111 </input>
<output>
<ID>OUT</ID>1132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>787</ID>
<type>AA_AND2</type>
<position>650.5,-96.5</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1113 </input>
<output>
<ID>OUT</ID>1133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>788</ID>
<type>AA_AND2</type>
<position>655.5,-93</position>
<input>
<ID>IN_0</ID>1116 </input>
<input>
<ID>IN_1</ID>1115 </input>
<output>
<ID>OUT</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>789</ID>
<type>AA_AND2</type>
<position>650.5,-89.5</position>
<input>
<ID>IN_0</ID>1118 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>790</ID>
<type>AA_AND2</type>
<position>655.5,-86</position>
<input>
<ID>IN_0</ID>1120 </input>
<input>
<ID>IN_1</ID>1119 </input>
<output>
<ID>OUT</ID>1136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>791</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-97.5</position>
<input>
<ID>IN_0</ID>1128 </input>
<input>
<ID>IN_1</ID>1136 </input>
<output>
<ID>OUT</ID>1144 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>792</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-102.5</position>
<input>
<ID>IN_0</ID>1127 </input>
<input>
<ID>IN_1</ID>1135 </input>
<output>
<ID>OUT</ID>1143 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>793</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-107.5</position>
<input>
<ID>IN_0</ID>1126 </input>
<input>
<ID>IN_1</ID>1134 </input>
<output>
<ID>OUT</ID>1142 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-112.5</position>
<input>
<ID>IN_0</ID>1125 </input>
<input>
<ID>IN_1</ID>1133 </input>
<output>
<ID>OUT</ID>1141 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>795</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-117.5</position>
<input>
<ID>IN_0</ID>1124 </input>
<input>
<ID>IN_1</ID>1132 </input>
<output>
<ID>OUT</ID>1140 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>796</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-122.5</position>
<input>
<ID>IN_0</ID>1123 </input>
<input>
<ID>IN_1</ID>1131 </input>
<output>
<ID>OUT</ID>1139 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>797</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-127.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<input>
<ID>IN_1</ID>1130 </input>
<output>
<ID>OUT</ID>1138 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>798</ID>
<type>AA_MUX_2x1</type>
<position>680.5,-132.5</position>
<input>
<ID>IN_0</ID>1121 </input>
<input>
<ID>IN_1</ID>1129 </input>
<output>
<ID>OUT</ID>1137 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>799</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>703,-114.5</position>
<input>
<ID>IN_0</ID>1137 </input>
<input>
<ID>IN_1</ID>1138 </input>
<input>
<ID>IN_2</ID>1139 </input>
<input>
<ID>IN_3</ID>1140 </input>
<input>
<ID>IN_4</ID>1141 </input>
<input>
<ID>IN_5</ID>1142 </input>
<input>
<ID>IN_6</ID>1143 </input>
<input>
<ID>IN_7</ID>1144 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_LABEL</type>
<position>680.5,-136</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>801</ID>
<type>AA_LABEL</type>
<position>681.5,-93.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>802</ID>
<type>GA_LED</type>
<position>694.5,-124.5</position>
<input>
<ID>N_in2</ID>1144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>803</ID>
<type>GA_LED</type>
<position>697,-124.5</position>
<input>
<ID>N_in2</ID>1143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>804</ID>
<type>GA_LED</type>
<position>699.5,-124.5</position>
<input>
<ID>N_in2</ID>1142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>805</ID>
<type>GA_LED</type>
<position>702,-124.5</position>
<input>
<ID>N_in2</ID>1141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>806</ID>
<type>GA_LED</type>
<position>704.5,-124.5</position>
<input>
<ID>N_in2</ID>1140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>807</ID>
<type>GA_LED</type>
<position>707,-124.5</position>
<input>
<ID>N_in2</ID>1139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>808</ID>
<type>GA_LED</type>
<position>709.5,-124.5</position>
<input>
<ID>N_in2</ID>1138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>809</ID>
<type>GA_LED</type>
<position>712,-124.5</position>
<input>
<ID>N_in2</ID>1137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>810</ID>
<type>AA_LABEL</type>
<position>712,-126.5</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>811</ID>
<type>AA_LABEL</type>
<position>709.5,-126.5</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>812</ID>
<type>AA_LABEL</type>
<position>707,-126.5</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>813</ID>
<type>AA_LABEL</type>
<position>704.5,-126.5</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>814</ID>
<type>AA_LABEL</type>
<position>702,-126.5</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>815</ID>
<type>AA_LABEL</type>
<position>699.5,-126.5</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>816</ID>
<type>AA_LABEL</type>
<position>697,-126.5</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>817</ID>
<type>AA_LABEL</type>
<position>694.5,-126.5</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>681</ID>
<type>AA_LABEL</type>
<position>625,-73</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>682</ID>
<type>AA_INVERTER</type>
<position>573,-38</position>
<input>
<ID>IN_0</ID>1082 </input>
<output>
<ID>OUT_0</ID>1083 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>683</ID>
<type>AA_TOGGLE</type>
<position>597.5,-13.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>684</ID>
<type>AA_LABEL</type>
<position>575,-45.5</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>685</ID>
<type>AA_LABEL</type>
<position>575,-47</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>686</ID>
<type>AE_REGISTER8</type>
<position>602,-29.5</position>
<input>
<ID>IN_0</ID>1020 </input>
<input>
<ID>IN_1</ID>1021 </input>
<input>
<ID>IN_2</ID>1022 </input>
<input>
<ID>IN_3</ID>1023 </input>
<input>
<ID>IN_4</ID>1024 </input>
<input>
<ID>IN_5</ID>1025 </input>
<input>
<ID>IN_6</ID>1026 </input>
<input>
<ID>IN_7</ID>1027 </input>
<output>
<ID>OUT_0</ID>1035 </output>
<output>
<ID>OUT_1</ID>1034 </output>
<output>
<ID>OUT_2</ID>1033 </output>
<output>
<ID>OUT_3</ID>1032 </output>
<output>
<ID>OUT_4</ID>1031 </output>
<output>
<ID>OUT_5</ID>1030 </output>
<output>
<ID>OUT_6</ID>1029 </output>
<output>
<ID>OUT_7</ID>1028 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1081 </input>
<input>
<ID>count_enable</ID>1043 </input>
<input>
<ID>count_up</ID>1043 </input>
<input>
<ID>load</ID>1083 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_REGISTER8</type>
<position>499,-89</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1152 </output>
<output>
<ID>OUT_1</ID>1151 </output>
<output>
<ID>OUT_2</ID>1150 </output>
<output>
<ID>OUT_3</ID>1149 </output>
<output>
<ID>OUT_4</ID>1148 </output>
<output>
<ID>OUT_5</ID>1147 </output>
<output>
<ID>OUT_6</ID>1146 </output>
<output>
<ID>OUT_7</ID>1145 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>1206 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>688</ID>
<type>AE_REGISTER8</type>
<position>619,-29.5</position>
<input>
<ID>IN_0</ID>1035 </input>
<input>
<ID>IN_1</ID>1034 </input>
<input>
<ID>IN_2</ID>1033 </input>
<input>
<ID>IN_3</ID>1032 </input>
<input>
<ID>IN_4</ID>1031 </input>
<input>
<ID>IN_5</ID>1030 </input>
<input>
<ID>IN_6</ID>1029 </input>
<input>
<ID>IN_7</ID>1028 </input>
<output>
<ID>OUT_0</ID>1046 </output>
<output>
<ID>OUT_1</ID>1045 </output>
<output>
<ID>OUT_2</ID>1041 </output>
<output>
<ID>OUT_3</ID>1040 </output>
<output>
<ID>OUT_4</ID>1039 </output>
<output>
<ID>OUT_5</ID>1038 </output>
<output>
<ID>OUT_6</ID>1037 </output>
<output>
<ID>OUT_7</ID>1036 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>1042 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_REGISTER8</type>
<position>499,-102</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1160 </output>
<output>
<ID>OUT_1</ID>1159 </output>
<output>
<ID>OUT_2</ID>1158 </output>
<output>
<ID>OUT_3</ID>1157 </output>
<output>
<ID>OUT_4</ID>1156 </output>
<output>
<ID>OUT_5</ID>1155 </output>
<output>
<ID>OUT_6</ID>1154 </output>
<output>
<ID>OUT_7</ID>1153 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>1207 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_REGISTER8</type>
<position>657,-68</position>
<input>
<ID>IN_0</ID>1070 </input>
<input>
<ID>IN_1</ID>1071 </input>
<input>
<ID>IN_2</ID>1072 </input>
<input>
<ID>IN_3</ID>1073 </input>
<input>
<ID>IN_4</ID>1074 </input>
<input>
<ID>IN_5</ID>1069 </input>
<input>
<ID>IN_6</ID>1076 </input>
<input>
<ID>IN_7</ID>1075 </input>
<output>
<ID>OUT_0</ID>1054 </output>
<output>
<ID>OUT_1</ID>1053 </output>
<output>
<ID>OUT_2</ID>1052 </output>
<output>
<ID>OUT_3</ID>1051 </output>
<output>
<ID>OUT_4</ID>1050 </output>
<output>
<ID>OUT_5</ID>1049 </output>
<output>
<ID>OUT_6</ID>1048 </output>
<output>
<ID>OUT_7</ID>1047 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>1044 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_RAM_8x8</type>
<position>634,-29</position>
<input>
<ID>ADDRESS_0</ID>1046 </input>
<input>
<ID>ADDRESS_1</ID>1045 </input>
<input>
<ID>ADDRESS_2</ID>1041 </input>
<input>
<ID>ADDRESS_3</ID>1040 </input>
<input>
<ID>ADDRESS_4</ID>1039 </input>
<input>
<ID>ADDRESS_5</ID>1038 </input>
<input>
<ID>ADDRESS_6</ID>1037 </input>
<input>
<ID>ADDRESS_7</ID>1036 </input>
<input>
<ID>DATA_IN_0</ID>1077 </input>
<input>
<ID>DATA_IN_1</ID>1062 </input>
<input>
<ID>DATA_IN_2</ID>1063 </input>
<input>
<ID>DATA_IN_3</ID>1064 </input>
<input>
<ID>DATA_IN_4</ID>1065 </input>
<input>
<ID>DATA_IN_5</ID>1066 </input>
<input>
<ID>DATA_IN_6</ID>1067 </input>
<input>
<ID>DATA_IN_7</ID>1068 </input>
<output>
<ID>DATA_OUT_0</ID>1077 </output>
<output>
<ID>DATA_OUT_1</ID>1062 </output>
<output>
<ID>DATA_OUT_2</ID>1063 </output>
<output>
<ID>DATA_OUT_3</ID>1064 </output>
<output>
<ID>DATA_OUT_4</ID>1065 </output>
<output>
<ID>DATA_OUT_5</ID>1066 </output>
<output>
<ID>DATA_OUT_6</ID>1067 </output>
<output>
<ID>DATA_OUT_7</ID>1068 </output>
<input>
<ID>ENABLE_0</ID>1061 </input>
<input>
<ID>write_enable</ID>1060 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_REGISTER8</type>
<position>674.5,-68</position>
<input>
<ID>IN_0</ID>1054 </input>
<input>
<ID>IN_1</ID>1053 </input>
<input>
<ID>IN_2</ID>1052 </input>
<input>
<ID>IN_3</ID>1051 </input>
<input>
<ID>IN_4</ID>1050 </input>
<input>
<ID>IN_5</ID>1049 </input>
<input>
<ID>IN_6</ID>1048 </input>
<input>
<ID>IN_7</ID>1047 </input>
<output>
<ID>OUT_0</ID>1056 </output>
<output>
<ID>OUT_1</ID>1057 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>1055 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>693</ID>
<type>DD_KEYPAD_HEX</type>
<position>582.5,-35.5</position>
<output>
<ID>OUT_0</ID>1020 </output>
<output>
<ID>OUT_1</ID>1021 </output>
<output>
<ID>OUT_2</ID>1022 </output>
<output>
<ID>OUT_3</ID>1023 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>694</ID>
<type>DD_KEYPAD_HEX</type>
<position>582.5,-23.5</position>
<output>
<ID>OUT_0</ID>1024 </output>
<output>
<ID>OUT_1</ID>1025 </output>
<output>
<ID>OUT_2</ID>1026 </output>
<output>
<ID>OUT_3</ID>1027 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>695</ID>
<type>BB_CLOCK</type>
<position>571,-61</position>
<output>
<ID>CLK</ID>1079 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>696</ID>
<type>AA_TOGGLE</type>
<position>600,-10.5</position>
<output>
<ID>OUT_0</ID>1043 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_LABEL</type>
<position>587.5,-12.5</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>698</ID>
<type>AA_LABEL</type>
<position>587.5,-10</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>699</ID>
<type>AA_TOGGLE</type>
<position>613,-13</position>
<output>
<ID>OUT_0</ID>1042 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>700</ID>
<type>AA_TOGGLE</type>
<position>601,-58</position>
<output>
<ID>OUT_0</ID>1059 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_LABEL</type>
<position>595.5,-55</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>702</ID>
<type>AA_TOGGLE</type>
<position>653.5,-60.5</position>
<output>
<ID>OUT_0</ID>1044 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>703</ID>
<type>AA_LABEL</type>
<position>597,-21.5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>704</ID>
<type>AA_LABEL</type>
<position>613.5,-21.5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>705</ID>
<type>AA_LABEL</type>
<position>634,-20.5</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>706</ID>
<type>AA_LABEL</type>
<position>657,-75.5</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>707</ID>
<type>AA_TOGGLE</type>
<position>671,-60.5</position>
<output>
<ID>OUT_0</ID>1055 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>626.5,-157.5</position>
<input>
<ID>IN_0</ID>831 </input>
<input>
<ID>IN_1</ID>762 </input>
<input>
<ID>IN_10</ID>765 </input>
<input>
<ID>IN_11</ID>757 </input>
<input>
<ID>IN_12</ID>764 </input>
<input>
<ID>IN_13</ID>756 </input>
<input>
<ID>IN_14</ID>763 </input>
<input>
<ID>IN_15</ID>755 </input>
<input>
<ID>IN_2</ID>830 </input>
<input>
<ID>IN_3</ID>761 </input>
<input>
<ID>IN_4</ID>768 </input>
<input>
<ID>IN_5</ID>760 </input>
<input>
<ID>IN_6</ID>767 </input>
<input>
<ID>IN_7</ID>759 </input>
<input>
<ID>IN_8</ID>766 </input>
<input>
<ID>IN_9</ID>758 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>708</ID>
<type>BE_ROM_8x8</type>
<position>687,-67.5</position>
<input>
<ID>ADDRESS_0</ID>1056 </input>
<input>
<ID>ADDRESS_1</ID>1057 </input>
<input>
<ID>ENABLE_0</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>130</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>626.5,-180.5</position>
<input>
<ID>IN_0</ID>831 </input>
<input>
<ID>IN_1</ID>762 </input>
<input>
<ID>IN_10</ID>765 </input>
<input>
<ID>IN_11</ID>757 </input>
<input>
<ID>IN_12</ID>764 </input>
<input>
<ID>IN_13</ID>756 </input>
<input>
<ID>IN_14</ID>763 </input>
<input>
<ID>IN_15</ID>755 </input>
<input>
<ID>IN_2</ID>830 </input>
<input>
<ID>IN_3</ID>761 </input>
<input>
<ID>IN_4</ID>768 </input>
<input>
<ID>IN_5</ID>760 </input>
<input>
<ID>IN_6</ID>767 </input>
<input>
<ID>IN_7</ID>759 </input>
<input>
<ID>IN_8</ID>766 </input>
<input>
<ID>IN_9</ID>758 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>709</ID>
<type>AA_TOGGLE</type>
<position>644,-26.5</position>
<output>
<ID>OUT_0</ID>1060 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_TOGGLE</type>
<position>644,-29.5</position>
<output>
<ID>OUT_0</ID>1061 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>586.5,-155.5</position>
<output>
<ID>OUT_0</ID>762 </output>
<output>
<ID>OUT_1</ID>761 </output>
<output>
<ID>OUT_2</ID>760 </output>
<output>
<ID>OUT_3</ID>759 </output>
<output>
<ID>OUT_4</ID>758 </output>
<output>
<ID>OUT_5</ID>757 </output>
<output>
<ID>OUT_6</ID>756 </output>
<output>
<ID>OUT_7</ID>755 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>711</ID>
<type>AA_LABEL</type>
<position>650.5,-26</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>712</ID>
<type>AA_LABEL</type>
<position>651,-29</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>586.5,-187</position>
<input>
<ID>ENABLE_0</ID>832 </input>
<output>
<ID>OUT_0</ID>831 </output>
<output>
<ID>OUT_1</ID>830 </output>
<output>
<ID>OUT_2</ID>768 </output>
<output>
<ID>OUT_3</ID>767 </output>
<output>
<ID>OUT_4</ID>766 </output>
<output>
<ID>OUT_5</ID>765 </output>
<output>
<ID>OUT_6</ID>764 </output>
<output>
<ID>OUT_7</ID>763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>713</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>647.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>1061 </input>
<input>
<ID>IN_0</ID>1077 </input>
<input>
<ID>IN_1</ID>1062 </input>
<input>
<ID>IN_2</ID>1063 </input>
<input>
<ID>IN_3</ID>1064 </input>
<input>
<ID>IN_4</ID>1065 </input>
<input>
<ID>IN_5</ID>1066 </input>
<input>
<ID>IN_6</ID>1067 </input>
<input>
<ID>IN_7</ID>1068 </input>
<output>
<ID>OUT_0</ID>1070 </output>
<output>
<ID>OUT_1</ID>1071 </output>
<output>
<ID>OUT_2</ID>1072 </output>
<output>
<ID>OUT_3</ID>1073 </output>
<output>
<ID>OUT_4</ID>1074 </output>
<output>
<ID>OUT_5</ID>1069 </output>
<output>
<ID>OUT_6</ID>1076 </output>
<output>
<ID>OUT_7</ID>1075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>714</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>625.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>1060 </input>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1175 </input>
<input>
<ID>IN_2</ID>1174 </input>
<input>
<ID>IN_3</ID>1173 </input>
<input>
<ID>IN_4</ID>1172 </input>
<input>
<ID>IN_5</ID>1171 </input>
<input>
<ID>IN_6</ID>1170 </input>
<input>
<ID>IN_7</ID>1169 </input>
<output>
<ID>OUT_0</ID>1077 </output>
<output>
<ID>OUT_1</ID>1062 </output>
<output>
<ID>OUT_2</ID>1063 </output>
<output>
<ID>OUT_3</ID>1064 </output>
<output>
<ID>OUT_4</ID>1065 </output>
<output>
<ID>OUT_5</ID>1066 </output>
<output>
<ID>OUT_6</ID>1067 </output>
<output>
<ID>OUT_7</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>136</ID>
<type>EE_VDD</type>
<position>586.5,-172</position>
<output>
<ID>OUT_0</ID>832 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>715</ID>
<type>AA_LABEL</type>
<position>674,-75.5</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>716</ID>
<type>AA_TOGGLE</type>
<position>696,-47</position>
<output>
<ID>OUT_0</ID>1078 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>717</ID>
<type>AA_LABEL</type>
<position>697.5,-44</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>718</ID>
<type>AA_AND2</type>
<position>597,-42.5</position>
<input>
<ID>IN_0</ID>1058 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>719</ID>
<type>AA_AND2</type>
<position>582.5,-60</position>
<input>
<ID>IN_0</ID>1080 </input>
<input>
<ID>IN_1</ID>1079 </input>
<output>
<ID>OUT</ID>1058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_TOGGLE</type>
<position>577,-57</position>
<output>
<ID>OUT_0</ID>1080 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>721</ID>
<type>AA_TOGGLE</type>
<position>568,-43.5</position>
<output>
<ID>OUT_0</ID>1082 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>722</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>637.5,-102</position>
<input>
<ID>ENABLE_0</ID>1087 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<output>
<ID>OUT_1</ID>1106 </output>
<output>
<ID>OUT_10</ID>1115 </output>
<output>
<ID>OUT_11</ID>1116 </output>
<output>
<ID>OUT_12</ID>1117 </output>
<output>
<ID>OUT_13</ID>1118 </output>
<output>
<ID>OUT_14</ID>1119 </output>
<output>
<ID>OUT_15</ID>1120 </output>
<output>
<ID>OUT_2</ID>1107 </output>
<output>
<ID>OUT_3</ID>1108 </output>
<output>
<ID>OUT_4</ID>1109 </output>
<output>
<ID>OUT_5</ID>1110 </output>
<output>
<ID>OUT_6</ID>1111 </output>
<output>
<ID>OUT_7</ID>1112 </output>
<output>
<ID>OUT_8</ID>1113 </output>
<output>
<ID>OUT_9</ID>1114 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>723</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>637.5,-125</position>
<input>
<ID>ENABLE_0</ID>1086 </input>
<output>
<ID>OUT_0</ID>1089 </output>
<output>
<ID>OUT_1</ID>1097 </output>
<output>
<ID>OUT_10</ID>1094 </output>
<output>
<ID>OUT_11</ID>1102 </output>
<output>
<ID>OUT_12</ID>1095 </output>
<output>
<ID>OUT_13</ID>1103 </output>
<output>
<ID>OUT_14</ID>1096 </output>
<output>
<ID>OUT_15</ID>1104 </output>
<output>
<ID>OUT_2</ID>1090 </output>
<output>
<ID>OUT_3</ID>1098 </output>
<output>
<ID>OUT_4</ID>1091 </output>
<output>
<ID>OUT_5</ID>1099 </output>
<output>
<ID>OUT_6</ID>1092 </output>
<output>
<ID>OUT_7</ID>1100 </output>
<output>
<ID>OUT_8</ID>1093 </output>
<output>
<ID>OUT_9</ID>1101 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>724</ID>
<type>AA_LABEL</type>
<position>598.5,-89</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>725</ID>
<type>AE_REGISTER8</type>
<position>499,-115.5</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1168 </output>
<output>
<ID>OUT_1</ID>1167 </output>
<output>
<ID>OUT_2</ID>1166 </output>
<output>
<ID>OUT_3</ID>1165 </output>
<output>
<ID>OUT_4</ID>1164 </output>
<output>
<ID>OUT_5</ID>1163 </output>
<output>
<ID>OUT_6</ID>1162 </output>
<output>
<ID>OUT_7</ID>1161 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>1208 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_REGISTER8</type>
<position>499,-128.5</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1184 </output>
<output>
<ID>OUT_1</ID>1175 </output>
<output>
<ID>OUT_2</ID>1174 </output>
<output>
<ID>OUT_3</ID>1173 </output>
<output>
<ID>OUT_4</ID>1172 </output>
<output>
<ID>OUT_5</ID>1171 </output>
<output>
<ID>OUT_6</ID>1170 </output>
<output>
<ID>OUT_7</ID>1169 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>1209 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-78</position>
<input>
<ID>IN_0</ID>1169 </input>
<input>
<ID>IN_1</ID>1161 </input>
<input>
<ID>IN_2</ID>1153 </input>
<input>
<ID>IN_3</ID>1145 </input>
<output>
<ID>OUT</ID>1176 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>728</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-89</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1162 </input>
<input>
<ID>IN_2</ID>1154 </input>
<input>
<ID>IN_3</ID>1146 </input>
<output>
<ID>OUT</ID>1177 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>729</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-100</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1163 </input>
<input>
<ID>IN_2</ID>1155 </input>
<input>
<ID>IN_3</ID>1147 </input>
<output>
<ID>OUT</ID>1178 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>730</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-109.5</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1164 </input>
<input>
<ID>IN_2</ID>1156 </input>
<input>
<ID>IN_3</ID>1148 </input>
<output>
<ID>OUT</ID>1179 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>731</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-120.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<input>
<ID>IN_1</ID>1165 </input>
<input>
<ID>IN_2</ID>1157 </input>
<input>
<ID>IN_3</ID>1149 </input>
<output>
<ID>OUT</ID>1180 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>732</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-131.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1166 </input>
<input>
<ID>IN_2</ID>1158 </input>
<input>
<ID>IN_3</ID>1150 </input>
<output>
<ID>OUT</ID>1181 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>733</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-142</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1167 </input>
<input>
<ID>IN_2</ID>1159 </input>
<input>
<ID>IN_3</ID>1151 </input>
<output>
<ID>OUT</ID>1182 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>734</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-153</position>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1168 </input>
<input>
<ID>IN_2</ID>1160 </input>
<input>
<ID>IN_3</ID>1152 </input>
<output>
<ID>OUT</ID>1183 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>735</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>563,-111</position>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1182 </input>
<input>
<ID>IN_2</ID>1181 </input>
<input>
<ID>IN_3</ID>1180 </input>
<input>
<ID>IN_4</ID>1179 </input>
<input>
<ID>IN_5</ID>1178 </input>
<input>
<ID>IN_6</ID>1177 </input>
<input>
<ID>IN_7</ID>1176 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>736</ID>
<type>DD_KEYPAD_HEX</type>
<position>466,-93</position>
<output>
<ID>OUT_0</ID>1186 </output>
<output>
<ID>OUT_1</ID>1187 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>737</ID>
<type>BB_CLOCK</type>
<position>487.5,-137</position>
<output>
<ID>CLK</ID>1185 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>738</ID>
<type>AA_LABEL</type>
<position>499.5,-121.5</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>739</ID>
<type>AA_LABEL</type>
<position>499.5,-108</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>740</ID>
<type>AA_LABEL</type>
<position>499.5,-95</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>741</ID>
<type>AA_LABEL</type>
<position>499.5,-81.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>742</ID>
<type>AA_LABEL</type>
<position>464.5,-86</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>743</ID>
<type>DD_KEYPAD_HEX</type>
<position>466,-107</position>
<output>
<ID>OUT_0</ID>1196 </output>
<output>
<ID>OUT_1</ID>1197 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>744</ID>
<type>AE_MUX_4x1</type>
<position>537,-78</position>
<input>
<ID>IN_0</ID>1169 </input>
<input>
<ID>IN_1</ID>1161 </input>
<input>
<ID>IN_2</ID>1153 </input>
<input>
<ID>IN_3</ID>1145 </input>
<output>
<ID>OUT</ID>1188 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>745</ID>
<type>AE_MUX_4x1</type>
<position>537,-89</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1162 </input>
<input>
<ID>IN_2</ID>1154 </input>
<input>
<ID>IN_3</ID>1146 </input>
<output>
<ID>OUT</ID>1189 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>746</ID>
<type>AE_MUX_4x1</type>
<position>537,-100</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1163 </input>
<input>
<ID>IN_2</ID>1155 </input>
<input>
<ID>IN_3</ID>1147 </input>
<output>
<ID>OUT</ID>1190 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>AE_MUX_4x1</type>
<position>537,-109.5</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1164 </input>
<input>
<ID>IN_2</ID>1156 </input>
<input>
<ID>IN_3</ID>1148 </input>
<output>
<ID>OUT</ID>1191 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>748</ID>
<type>AE_MUX_4x1</type>
<position>537,-120.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<input>
<ID>IN_1</ID>1165 </input>
<input>
<ID>IN_2</ID>1157 </input>
<input>
<ID>IN_3</ID>1149 </input>
<output>
<ID>OUT</ID>1192 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>749</ID>
<type>AE_MUX_4x1</type>
<position>537,-131.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1166 </input>
<input>
<ID>IN_2</ID>1158 </input>
<input>
<ID>IN_3</ID>1150 </input>
<output>
<ID>OUT</ID>1193 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>750</ID>
<type>AE_MUX_4x1</type>
<position>537,-142</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1167 </input>
<input>
<ID>IN_2</ID>1159 </input>
<input>
<ID>IN_3</ID>1151 </input>
<output>
<ID>OUT</ID>1194 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_MUX_4x1</type>
<position>537,-153</position>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1168 </input>
<input>
<ID>IN_2</ID>1160 </input>
<input>
<ID>IN_3</ID>1152 </input>
<output>
<ID>OUT</ID>1195 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>752</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>565,-121.5</position>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1194 </input>
<input>
<ID>IN_2</ID>1193 </input>
<input>
<ID>IN_3</ID>1192 </input>
<input>
<ID>IN_4</ID>1191 </input>
<input>
<ID>IN_5</ID>1190 </input>
<input>
<ID>IN_6</ID>1189 </input>
<input>
<ID>IN_7</ID>1188 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 36</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>753</ID>
<type>AA_LABEL</type>
<position>464.5,-100</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>754</ID>
<type>DD_KEYPAD_HEX</type>
<position>482,-106.5</position>
<output>
<ID>OUT_0</ID>1201 </output>
<output>
<ID>OUT_1</ID>1200 </output>
<output>
<ID>OUT_2</ID>1199 </output>
<output>
<ID>OUT_3</ID>1198 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>755</ID>
<type>DD_KEYPAD_HEX</type>
<position>482,-118.5</position>
<output>
<ID>OUT_0</ID>1205 </output>
<output>
<ID>OUT_1</ID>1204 </output>
<output>
<ID>OUT_2</ID>1203 </output>
<output>
<ID>OUT_3</ID>1202 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>756</ID>
<type>AA_LABEL</type>
<position>482,-99.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>757</ID>
<type>BA_DECODER_2x4</type>
<position>484,-73.5</position>
<input>
<ID>ENABLE</ID>1210 </input>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT_0</ID>1206 </output>
<output>
<ID>OUT_1</ID>1207 </output>
<output>
<ID>OUT_2</ID>1208 </output>
<output>
<ID>OUT_3</ID>1209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>AA_TOGGLE</type>
<position>478,-73</position>
<output>
<ID>OUT_0</ID>1210 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>759</ID>
<type>AA_LABEL</type>
<position>475.5,-72.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>760</ID>
<type>DD_KEYPAD_HEX</type>
<position>479,-86</position>
<output>
<ID>OUT_0</ID>196 </output>
<output>
<ID>OUT_1</ID>195 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_LABEL</type>
<position>479.5,-79</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>762</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>581,-100</position>
<input>
<ID>ENABLE_0</ID>1213 </input>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1182 </input>
<input>
<ID>IN_2</ID>1181 </input>
<input>
<ID>IN_3</ID>1180 </input>
<input>
<ID>IN_4</ID>1179 </input>
<input>
<ID>IN_5</ID>1178 </input>
<input>
<ID>IN_6</ID>1177 </input>
<input>
<ID>IN_7</ID>1176 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>763</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>581,-131.5</position>
<input>
<ID>ENABLE_0</ID>1214 </input>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1194 </input>
<input>
<ID>IN_2</ID>1193 </input>
<input>
<ID>IN_3</ID>1192 </input>
<input>
<ID>IN_4</ID>1191 </input>
<input>
<ID>IN_5</ID>1190 </input>
<input>
<ID>IN_6</ID>1189 </input>
<input>
<ID>IN_7</ID>1188 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>764</ID>
<type>EE_VDD</type>
<position>581,-88</position>
<output>
<ID>OUT_0</ID>1213 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_LABEL</type>
<position>578.5,-91</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>766</ID>
<type>AA_LABEL</type>
<position>556,-104.5</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>767</ID>
<type>AA_LABEL</type>
<position>581,-137.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>768</ID>
<type>AA_LABEL</type>
<position>556,-115.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>769</ID>
<type>EE_VDD</type>
<position>581,-116.5</position>
<output>
<ID>OUT_0</ID>1214 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>770</ID>
<type>BA_DECODER_2x4</type>
<position>629,-85.5</position>
<input>
<ID>ENABLE</ID>1084 </input>
<input>
<ID>IN_0</ID>1085 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<output>
<ID>OUT_1</ID>1087 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>AA_TOGGLE</type>
<position>624,-84</position>
<output>
<ID>OUT_0</ID>1084 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515.5,-143,515.5,-117.5</points>
<intersection>-143 1</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,-143,534,-143</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<intersection>515.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-117.5,515.5,-117.5</points>
<connection>
<GID>725</GID>
<name>OUT_1</name></connection>
<intersection>515.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516,-154,516,-118.5</points>
<intersection>-154 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,-118.5,516,-118.5</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>516 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>516,-154,534,-154</points>
<connection>
<GID>734</GID>
<name>IN_1</name></connection>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<intersection>516 0</intersection></hsegment></shape></wire>
<wire>
<ID>1169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517.5,-162,517.5,-124.5</points>
<intersection>-162 1</intersection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517.5,-162,572,-162</points>
<intersection>517.5 0</intersection>
<intersection>521.5 5</intersection>
<intersection>572 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-124.5,517.5,-124.5</points>
<connection>
<GID>726</GID>
<name>OUT_7</name></connection>
<intersection>517.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>572,-162,572,-64</points>
<intersection>-162 1</intersection>
<intersection>-64 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>521.5,-162,521.5,-81</points>
<intersection>-162 1</intersection>
<intersection>-81 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>572,-64,623.5,-64</points>
<connection>
<GID>714</GID>
<name>IN_7</name></connection>
<intersection>572 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>521.5,-81,534,-81</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>521.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518,-161.5,518,-125.5</points>
<intersection>-161.5 1</intersection>
<intersection>-125.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>518,-161.5,572.5,-161.5</points>
<intersection>518 0</intersection>
<intersection>521.5 7</intersection>
<intersection>572.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-125.5,518,-125.5</points>
<connection>
<GID>726</GID>
<name>OUT_6</name></connection>
<intersection>518 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>572.5,-161.5,572.5,-65</points>
<intersection>-161.5 1</intersection>
<intersection>-65 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>572.5,-65,623.5,-65</points>
<connection>
<GID>714</GID>
<name>IN_6</name></connection>
<intersection>572.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>521.5,-161.5,521.5,-92</points>
<intersection>-161.5 1</intersection>
<intersection>-92 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>521.5,-92,534,-92</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>521.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>518.5,-161,518.5,-126.5</points>
<intersection>-161 1</intersection>
<intersection>-126.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>518.5,-161,573,-161</points>
<intersection>518.5 0</intersection>
<intersection>521.5 8</intersection>
<intersection>573 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-126.5,518.5,-126.5</points>
<connection>
<GID>726</GID>
<name>OUT_5</name></connection>
<intersection>518.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>573,-161,573,-66</points>
<intersection>-161 1</intersection>
<intersection>-66 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>573,-66,623.5,-66</points>
<connection>
<GID>714</GID>
<name>IN_5</name></connection>
<intersection>573 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>521.5,-161,521.5,-103</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>-161 1</intersection>
<intersection>-103 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>521.5,-103,534,-103</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>521.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-160.5,573.5,-160.5</points>
<intersection>519 6</intersection>
<intersection>521.5 13</intersection>
<intersection>573.5 11</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>519,-160.5,519,-127.5</points>
<intersection>-160.5 1</intersection>
<intersection>-127.5 15</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>573.5,-160.5,573.5,-67</points>
<intersection>-160.5 1</intersection>
<intersection>-67 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>573.5,-67,623.5,-67</points>
<connection>
<GID>714</GID>
<name>IN_4</name></connection>
<intersection>573.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>521.5,-160.5,521.5,-112.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection>
<intersection>-112.5 16</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>503,-127.5,519,-127.5</points>
<connection>
<GID>726</GID>
<name>OUT_4</name></connection>
<intersection>519 6</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>521.5,-112.5,534,-112.5</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>521.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>1173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521,-158.5,521,-123.5</points>
<intersection>-158.5 1</intersection>
<intersection>-128.5 2</intersection>
<intersection>-123.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>521,-158.5,574,-158.5</points>
<intersection>521 0</intersection>
<intersection>521.5 10</intersection>
<intersection>574 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-128.5,521,-128.5</points>
<connection>
<GID>726</GID>
<name>OUT_3</name></connection>
<intersection>521 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>574,-158.5,574,-68</points>
<intersection>-158.5 1</intersection>
<intersection>-68 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>574,-68,623.5,-68</points>
<connection>
<GID>714</GID>
<name>IN_3</name></connection>
<intersection>574 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>521.5,-158.5,521.5,-123.5</points>
<intersection>-158.5 1</intersection>
<intersection>-123.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>521,-123.5,534,-123.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>521 0</intersection>
<intersection>521.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>1174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>519.5,-160,519.5,-129.5</points>
<intersection>-160 1</intersection>
<intersection>-129.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>519.5,-160,574.5,-160</points>
<intersection>519.5 0</intersection>
<intersection>521.5 4</intersection>
<intersection>574.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-129.5,519.5,-129.5</points>
<connection>
<GID>726</GID>
<name>OUT_2</name></connection>
<intersection>519.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>574.5,-160,574.5,-69</points>
<intersection>-160 1</intersection>
<intersection>-69 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>521.5,-160,521.5,-134.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<intersection>-160 1</intersection>
<intersection>-134.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>574.5,-69,623.5,-69</points>
<connection>
<GID>714</GID>
<name>IN_2</name></connection>
<intersection>574.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>521.5,-134.5,534,-134.5</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>521.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520,-159.5,520,-130.5</points>
<intersection>-159.5 1</intersection>
<intersection>-130.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520,-159.5,575,-159.5</points>
<intersection>520 0</intersection>
<intersection>521.5 8</intersection>
<intersection>575 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-130.5,520,-130.5</points>
<connection>
<GID>726</GID>
<name>OUT_1</name></connection>
<intersection>520 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>575,-159.5,575,-70</points>
<intersection>-159.5 1</intersection>
<intersection>-70 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>575,-70,623.5,-70</points>
<connection>
<GID>714</GID>
<name>IN_1</name></connection>
<intersection>575 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>521.5,-159.5,521.5,-145</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>-159.5 1</intersection>
<intersection>-145 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>521.5,-145,534,-145</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>521.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-107,546,-78</points>
<intersection>-107 2</intersection>
<intersection>-96.5 3</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-78,546,-78</points>
<connection>
<GID>727</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-107,558,-107</points>
<connection>
<GID>735</GID>
<name>IN_7</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>546,-96.5,579,-96.5</points>
<connection>
<GID>762</GID>
<name>IN_7</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>1177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-108,546,-89</points>
<intersection>-108 2</intersection>
<intersection>-97.5 4</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-89,546,-89</points>
<connection>
<GID>728</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-108,558,-108</points>
<connection>
<GID>735</GID>
<name>IN_6</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>546,-97.5,579,-97.5</points>
<connection>
<GID>762</GID>
<name>IN_6</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>1178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-109,546,-98.5</points>
<intersection>-109 2</intersection>
<intersection>-100 1</intersection>
<intersection>-98.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-100,546,-100</points>
<connection>
<GID>729</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-109,558,-109</points>
<connection>
<GID>735</GID>
<name>IN_5</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>546,-98.5,579,-98.5</points>
<connection>
<GID>762</GID>
<name>IN_5</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>1179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-109.5,558,-109.5</points>
<connection>
<GID>730</GID>
<name>OUT</name></connection>
<intersection>547 4</intersection>
<intersection>558 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>547,-109.5,547,-99.5</points>
<intersection>-109.5 1</intersection>
<intersection>-99.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>547,-99.5,579,-99.5</points>
<connection>
<GID>762</GID>
<name>IN_4</name></connection>
<intersection>547 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>558,-110,558,-109.5</points>
<connection>
<GID>735</GID>
<name>IN_4</name></connection>
<intersection>-109.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-120.5,546,-111</points>
<intersection>-120.5 1</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-120.5,546,-120.5</points>
<connection>
<GID>731</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-111,558,-111</points>
<connection>
<GID>735</GID>
<name>IN_3</name></connection>
<intersection>546 0</intersection>
<intersection>548 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>548,-111,548,-100.5</points>
<intersection>-111 2</intersection>
<intersection>-100.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>548,-100.5,579,-100.5</points>
<connection>
<GID>762</GID>
<name>IN_3</name></connection>
<intersection>548 3</intersection></hsegment></shape></wire>
<wire>
<ID>1181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-131.5,546,-112</points>
<intersection>-131.5 1</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-131.5,546,-131.5</points>
<connection>
<GID>732</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-112,558,-112</points>
<connection>
<GID>735</GID>
<name>IN_2</name></connection>
<intersection>546 0</intersection>
<intersection>549 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>549,-112,549,-101.5</points>
<intersection>-112 2</intersection>
<intersection>-101.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>549,-101.5,579,-101.5</points>
<connection>
<GID>762</GID>
<name>IN_2</name></connection>
<intersection>549 3</intersection></hsegment></shape></wire>
<wire>
<ID>1182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-142,546,-113</points>
<intersection>-142 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-142,546,-142</points>
<connection>
<GID>733</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-113,558,-113</points>
<connection>
<GID>735</GID>
<name>IN_1</name></connection>
<intersection>546 0</intersection>
<intersection>550 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>550,-113,550,-102.5</points>
<intersection>-113 2</intersection>
<intersection>-102.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>550,-102.5,579,-102.5</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>550 3</intersection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-153,546,-114</points>
<intersection>-153 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>546,-114,558,-114</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>546 0</intersection>
<intersection>551 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527.5,-153,546,-153</points>
<connection>
<GID>734</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>551,-114,551,-103.5</points>
<intersection>-114 1</intersection>
<intersection>-103.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>551,-103.5,579,-103.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>551 3</intersection></hsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-159,520.5,-131.5</points>
<intersection>-159 1</intersection>
<intersection>-131.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520.5,-159,575.5,-159</points>
<intersection>520.5 0</intersection>
<intersection>521.5 14</intersection>
<intersection>575.5 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-131.5,520.5,-131.5</points>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection>
<intersection>520.5 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>575.5,-159,575.5,-71</points>
<intersection>-159 1</intersection>
<intersection>-71 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>521.5,-159,521.5,-156</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection>
<intersection>-156 17</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>575.5,-71,623.5,-71</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>575.5 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>521.5,-156,534,-156</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>521.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>494.5,-137,494.5,-94</points>
<intersection>-137 10</intersection>
<intersection>-133.5 8</intersection>
<intersection>-120.5 7</intersection>
<intersection>-107 6</intersection>
<intersection>-94 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>494.5,-94,498,-94</points>
<connection>
<GID>687</GID>
<name>clock</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>494.5,-107,498,-107</points>
<connection>
<GID>689</GID>
<name>clock</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>494.5,-120.5,498,-120.5</points>
<connection>
<GID>725</GID>
<name>clock</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>494.5,-133.5,498,-133.5</points>
<connection>
<GID>726</GID>
<name>clock</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>491.5,-137,494.5,-137</points>
<connection>
<GID>737</GID>
<name>CLK</name></connection>
<intersection>494.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525.5,-148,525.5,-70</points>
<connection>
<GID>734</GID>
<name>SEL_0</name></connection>
<connection>
<GID>733</GID>
<name>SEL_0</name></connection>
<connection>
<GID>732</GID>
<name>SEL_0</name></connection>
<connection>
<GID>731</GID>
<name>SEL_0</name></connection>
<connection>
<GID>730</GID>
<name>SEL_0</name></connection>
<connection>
<GID>729</GID>
<name>SEL_0</name></connection>
<connection>
<GID>728</GID>
<name>SEL_0</name></connection>
<connection>
<GID>727</GID>
<name>SEL_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>472,-70,525.5,-70</points>
<intersection>472 2</intersection>
<intersection>525.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>472,-96,472,-70</points>
<intersection>-96 3</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>471,-96,472,-96</points>
<connection>
<GID>736</GID>
<name>OUT_0</name></connection>
<intersection>472 2</intersection></hsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,-148,524.5,-69.5</points>
<connection>
<GID>734</GID>
<name>SEL_1</name></connection>
<connection>
<GID>733</GID>
<name>SEL_1</name></connection>
<connection>
<GID>732</GID>
<name>SEL_1</name></connection>
<connection>
<GID>731</GID>
<name>SEL_1</name></connection>
<connection>
<GID>730</GID>
<name>SEL_1</name></connection>
<connection>
<GID>729</GID>
<name>SEL_1</name></connection>
<connection>
<GID>728</GID>
<name>SEL_1</name></connection>
<connection>
<GID>727</GID>
<name>SEL_1</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>471.5,-69.5,524.5,-69.5</points>
<intersection>471.5 2</intersection>
<intersection>524.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>471.5,-94,471.5,-69.5</points>
<intersection>-94 3</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>471,-94,471.5,-94</points>
<connection>
<GID>736</GID>
<name>OUT_1</name></connection>
<intersection>471.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-117.5,540.5,-78</points>
<intersection>-117.5 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-78,540.5,-78</points>
<connection>
<GID>744</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-117.5,560,-117.5</points>
<connection>
<GID>752</GID>
<name>IN_7</name></connection>
<intersection>540.5 0</intersection>
<intersection>546.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>546.5,-128,546.5,-117.5</points>
<intersection>-128 4</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>546.5,-128,579,-128</points>
<connection>
<GID>763</GID>
<name>IN_7</name></connection>
<intersection>546.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-118.5,540.5,-89</points>
<intersection>-118.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-89,540.5,-89</points>
<connection>
<GID>745</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-118.5,560,-118.5</points>
<connection>
<GID>752</GID>
<name>IN_6</name></connection>
<intersection>540.5 0</intersection>
<intersection>547 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>547,-129,547,-118.5</points>
<intersection>-129 4</intersection>
<intersection>-118.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>547,-129,579,-129</points>
<connection>
<GID>763</GID>
<name>IN_6</name></connection>
<intersection>547 3</intersection></hsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-119.5,540.5,-100</points>
<intersection>-119.5 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-100,540.5,-100</points>
<connection>
<GID>746</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-119.5,560,-119.5</points>
<connection>
<GID>752</GID>
<name>IN_5</name></connection>
<intersection>540.5 0</intersection>
<intersection>549 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>549,-130,549,-119.5</points>
<intersection>-130 4</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>549,-130,579,-130</points>
<connection>
<GID>763</GID>
<name>IN_5</name></connection>
<intersection>549 3</intersection></hsegment></shape></wire>
<wire>
<ID>1191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-120.5,540.5,-109.5</points>
<intersection>-120.5 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-109.5,540.5,-109.5</points>
<connection>
<GID>747</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-120.5,560,-120.5</points>
<connection>
<GID>752</GID>
<name>IN_4</name></connection>
<intersection>540.5 0</intersection>
<intersection>550.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>550.5,-131,550.5,-120.5</points>
<intersection>-131 4</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>550.5,-131,579,-131</points>
<connection>
<GID>763</GID>
<name>IN_4</name></connection>
<intersection>550.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>540.5,-121.5,560,-121.5</points>
<connection>
<GID>752</GID>
<name>IN_3</name></connection>
<intersection>540.5 2</intersection>
<intersection>552.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>540.5,-121.5,540.5,-120.5</points>
<intersection>-121.5 1</intersection>
<intersection>-120.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>540,-120.5,540.5,-120.5</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<intersection>540.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>552.5,-132,552.5,-121.5</points>
<intersection>-132 5</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>552.5,-132,579,-132</points>
<connection>
<GID>763</GID>
<name>IN_3</name></connection>
<intersection>552.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-131.5,540.5,-122.5</points>
<intersection>-131.5 1</intersection>
<intersection>-122.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-131.5,540.5,-131.5</points>
<connection>
<GID>749</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-122.5,560,-122.5</points>
<connection>
<GID>752</GID>
<name>IN_2</name></connection>
<intersection>540.5 0</intersection>
<intersection>554.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>554.5,-133,554.5,-122.5</points>
<intersection>-133 4</intersection>
<intersection>-122.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>554.5,-133,579,-133</points>
<connection>
<GID>763</GID>
<name>IN_2</name></connection>
<intersection>554.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-142,540.5,-123.5</points>
<intersection>-142 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-142,540.5,-142</points>
<connection>
<GID>750</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-123.5,560,-123.5</points>
<connection>
<GID>752</GID>
<name>IN_1</name></connection>
<intersection>540.5 0</intersection>
<intersection>555.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>555.5,-134,555.5,-123.5</points>
<intersection>-134 4</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>555.5,-134,579,-134</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<intersection>555.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-153,540.5,-124.5</points>
<intersection>-153 2</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540.5,-124.5,560,-124.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection>
<intersection>556.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540,-153,540.5,-153</points>
<connection>
<GID>751</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>556.5,-135,556.5,-124.5</points>
<intersection>-135 4</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>556.5,-135,579,-135</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>556.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538,-148,538,-71</points>
<connection>
<GID>751</GID>
<name>SEL_0</name></connection>
<connection>
<GID>750</GID>
<name>SEL_0</name></connection>
<connection>
<GID>749</GID>
<name>SEL_0</name></connection>
<connection>
<GID>748</GID>
<name>SEL_0</name></connection>
<connection>
<GID>747</GID>
<name>SEL_0</name></connection>
<connection>
<GID>746</GID>
<name>SEL_0</name></connection>
<connection>
<GID>745</GID>
<name>SEL_0</name></connection>
<connection>
<GID>744</GID>
<name>SEL_0</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>473,-71,538,-71</points>
<intersection>473 2</intersection>
<intersection>538 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>473,-110,473,-71</points>
<intersection>-110 3</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>471,-110,473,-110</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>473 2</intersection></hsegment></shape></wire>
<wire>
<ID>1197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,-148,537,-70.5</points>
<connection>
<GID>751</GID>
<name>SEL_1</name></connection>
<connection>
<GID>750</GID>
<name>SEL_1</name></connection>
<connection>
<GID>749</GID>
<name>SEL_1</name></connection>
<connection>
<GID>748</GID>
<name>SEL_1</name></connection>
<connection>
<GID>747</GID>
<name>SEL_1</name></connection>
<connection>
<GID>746</GID>
<name>SEL_1</name></connection>
<connection>
<GID>745</GID>
<name>SEL_1</name></connection>
<connection>
<GID>744</GID>
<name>SEL_1</name></connection>
<intersection>-70.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>472.5,-70.5,537,-70.5</points>
<intersection>472.5 16</intersection>
<intersection>537 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>472.5,-108,472.5,-70.5</points>
<intersection>-108 18</intersection>
<intersection>-70.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>471,-108,472.5,-108</points>
<connection>
<GID>743</GID>
<name>OUT_1</name></connection>
<intersection>472.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>1198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-124.5,493.5,-85</points>
<intersection>-124.5 6</intersection>
<intersection>-111.5 3</intersection>
<intersection>-103.5 4</intersection>
<intersection>-98 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493.5,-85,495,-85</points>
<connection>
<GID>687</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>493.5,-98,495,-98</points>
<connection>
<GID>689</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>493.5,-111.5,495,-111.5</points>
<connection>
<GID>725</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>487,-103.5,493.5,-103.5</points>
<connection>
<GID>754</GID>
<name>OUT_3</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>493.5,-124.5,495,-124.5</points>
<connection>
<GID>726</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,-125.5,493,-86</points>
<intersection>-125.5 6</intersection>
<intersection>-112.5 5</intersection>
<intersection>-105.5 2</intersection>
<intersection>-99 3</intersection>
<intersection>-86 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>487,-105.5,493,-105.5</points>
<connection>
<GID>754</GID>
<name>OUT_2</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>493,-99,495,-99</points>
<connection>
<GID>689</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>493,-86,495,-86</points>
<connection>
<GID>687</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>493,-112.5,495,-112.5</points>
<connection>
<GID>725</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>493,-125.5,495,-125.5</points>
<connection>
<GID>726</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment></shape></wire>
<wire>
<ID>1200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,-126.5,492.5,-87</points>
<intersection>-126.5 6</intersection>
<intersection>-113.5 3</intersection>
<intersection>-107.5 2</intersection>
<intersection>-100 4</intersection>
<intersection>-87 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>487,-107.5,492.5,-107.5</points>
<connection>
<GID>754</GID>
<name>OUT_1</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>492.5,-113.5,495,-113.5</points>
<connection>
<GID>725</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>492.5,-100,495,-100</points>
<connection>
<GID>689</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>492.5,-87,495,-87</points>
<connection>
<GID>687</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>492.5,-126.5,495,-126.5</points>
<connection>
<GID>726</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492,-127.5,492,-88</points>
<intersection>-127.5 6</intersection>
<intersection>-114.5 3</intersection>
<intersection>-109.5 2</intersection>
<intersection>-101 4</intersection>
<intersection>-88 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>487,-109.5,492,-109.5</points>
<connection>
<GID>754</GID>
<name>OUT_0</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>492,-114.5,495,-114.5</points>
<connection>
<GID>725</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>492,-101,495,-101</points>
<connection>
<GID>689</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>492,-88,495,-88</points>
<connection>
<GID>687</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>492,-127.5,495,-127.5</points>
<connection>
<GID>726</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,-128.5,491.5,-89</points>
<intersection>-128.5 5</intersection>
<intersection>-115.5 2</intersection>
<intersection>-102 3</intersection>
<intersection>-89 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>487,-115.5,495,-115.5</points>
<connection>
<GID>725</GID>
<name>IN_3</name></connection>
<connection>
<GID>755</GID>
<name>OUT_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>491.5,-102,495,-102</points>
<connection>
<GID>689</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>491.5,-89,495,-89</points>
<connection>
<GID>687</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491.5,-128.5,495,-128.5</points>
<connection>
<GID>726</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,-129.5,491,-90</points>
<intersection>-129.5 5</intersection>
<intersection>-117.5 2</intersection>
<intersection>-116.5 4</intersection>
<intersection>-103 3</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,-90,495,-90</points>
<connection>
<GID>687</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>487,-117.5,491,-117.5</points>
<connection>
<GID>755</GID>
<name>OUT_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>491,-103,495,-103</points>
<connection>
<GID>689</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>491,-116.5,495,-116.5</points>
<connection>
<GID>725</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491,-129.5,495,-129.5</points>
<connection>
<GID>726</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490.5,-130.5,490.5,-91</points>
<intersection>-130.5 5</intersection>
<intersection>-119.5 2</intersection>
<intersection>-117.5 4</intersection>
<intersection>-104 3</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>490.5,-91,495,-91</points>
<connection>
<GID>687</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>487,-119.5,490.5,-119.5</points>
<connection>
<GID>755</GID>
<name>OUT_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>490.5,-104,495,-104</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490.5,-117.5,495,-117.5</points>
<connection>
<GID>725</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>490.5,-130.5,495,-130.5</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490,-131.5,490,-92</points>
<intersection>-131.5 5</intersection>
<intersection>-121.5 2</intersection>
<intersection>-118.5 4</intersection>
<intersection>-105 3</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>490,-92,495,-92</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>487,-121.5,490,-121.5</points>
<connection>
<GID>755</GID>
<name>OUT_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>490,-105,495,-105</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490,-118.5,495,-118.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>490,-131.5,495,-131.5</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-83,497,-75</points>
<intersection>-83 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-75,497,-75</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-83,498,-83</points>
<connection>
<GID>687</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-96,497,-74</points>
<intersection>-96 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-74,497,-74</points>
<connection>
<GID>757</GID>
<name>OUT_1</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-96,498,-96</points>
<connection>
<GID>689</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-109.5,497,-73</points>
<intersection>-109.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-73,497,-73</points>
<connection>
<GID>757</GID>
<name>OUT_2</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-109.5,498,-109.5</points>
<connection>
<GID>725</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-122.5,497,-72</points>
<intersection>-122.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-72,497,-72</points>
<connection>
<GID>757</GID>
<name>OUT_3</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-122.5,498,-122.5</points>
<connection>
<GID>726</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>480,-73,481,-73</points>
<connection>
<GID>758</GID>
<name>OUT_0</name></connection>
<intersection>481 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>481,-73,481,-72</points>
<connection>
<GID>757</GID>
<name>ENABLE</name></connection>
<intersection>-73 1</intersection></vsegment></shape></wire>
<wire>
<ID>1213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,-95,581,-89</points>
<connection>
<GID>764</GID>
<name>OUT_0</name></connection>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,-126.5,581,-117.5</points>
<connection>
<GID>769</GID>
<name>OUT_0</name></connection>
<connection>
<GID>763</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-189.5,592.5,-186</points>
<intersection>-189.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-186,624.5,-186</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>592.5 0</intersection>
<intersection>606 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-189.5,592.5,-189.5</points>
<connection>
<GID>134</GID>
<name>OUT_1</name></connection>
<intersection>592.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>606,-186,606,-163</points>
<intersection>-186 1</intersection>
<intersection>-163 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>606,-163,624.5,-163</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>606 3</intersection></hsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,-190.5,593,-188</points>
<intersection>-190.5 2</intersection>
<intersection>-188 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>593,-188,624.5,-188</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>593 0</intersection>
<intersection>607 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-190.5,593,-190.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>593 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>607,-188,607,-165</points>
<intersection>-188 1</intersection>
<intersection>-165 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>607,-165,624.5,-165</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>607 3</intersection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586.5,-182,586.5,-173</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<connection>
<GID>134</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485.5,-87,485.5,-78.5</points>
<intersection>-87 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,-87,485.5,-87</points>
<connection>
<GID>760</GID>
<name>OUT_1</name></connection>
<intersection>485.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>478.5,-78.5,485.5,-78.5</points>
<intersection>478.5 3</intersection>
<intersection>485.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>478.5,-78.5,478.5,-75</points>
<intersection>-78.5 2</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>478.5,-75,481,-75</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>478.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487.5,-89,487.5,-76.5</points>
<intersection>-89 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,-89,487.5,-89</points>
<connection>
<GID>760</GID>
<name>OUT_0</name></connection>
<intersection>487.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>480.5,-76.5,487.5,-76.5</points>
<intersection>480.5 3</intersection>
<intersection>487.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>480.5,-76.5,480.5,-74</points>
<intersection>-76.5 2</intersection>
<intersection>-74 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>480.5,-74,481,-74</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<intersection>480.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-38.5,592.5,-32.5</points>
<intersection>-38.5 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-32.5,598,-32.5</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-38.5,592.5,-38.5</points>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-36.5,592.5,-31.5</points>
<intersection>-36.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-31.5,598,-31.5</points>
<connection>
<GID>686</GID>
<name>IN_1</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-36.5,592.5,-36.5</points>
<connection>
<GID>693</GID>
<name>OUT_1</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-34.5,592.5,-30.5</points>
<intersection>-34.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-30.5,598,-30.5</points>
<connection>
<GID>686</GID>
<name>IN_2</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-34.5,592.5,-34.5</points>
<connection>
<GID>693</GID>
<name>OUT_2</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-32.5,592.5,-29.5</points>
<intersection>-32.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-29.5,598,-29.5</points>
<connection>
<GID>686</GID>
<name>IN_3</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-32.5,592.5,-32.5</points>
<connection>
<GID>693</GID>
<name>OUT_3</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-28.5,592.5,-26.5</points>
<intersection>-28.5 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-28.5,598,-28.5</points>
<connection>
<GID>686</GID>
<name>IN_4</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-26.5,592.5,-26.5</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-27.5,592.5,-24.5</points>
<intersection>-27.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-27.5,598,-27.5</points>
<connection>
<GID>686</GID>
<name>IN_5</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-24.5,592.5,-24.5</points>
<connection>
<GID>694</GID>
<name>OUT_1</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-26.5,592.5,-22.5</points>
<intersection>-26.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-26.5,598,-26.5</points>
<connection>
<GID>686</GID>
<name>IN_6</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>587.5,-22.5,592.5,-22.5</points>
<connection>
<GID>694</GID>
<name>OUT_2</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>587.5,-25.5,598,-25.5</points>
<connection>
<GID>686</GID>
<name>IN_7</name></connection>
<intersection>587.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>587.5,-25.5,587.5,-20.5</points>
<connection>
<GID>694</GID>
<name>OUT_3</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-25.5,615,-25.5</points>
<connection>
<GID>686</GID>
<name>OUT_7</name></connection>
<connection>
<GID>688</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-26.5,615,-26.5</points>
<connection>
<GID>686</GID>
<name>OUT_6</name></connection>
<connection>
<GID>688</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-27.5,615,-27.5</points>
<connection>
<GID>686</GID>
<name>OUT_5</name></connection>
<connection>
<GID>688</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-28.5,615,-28.5</points>
<connection>
<GID>686</GID>
<name>OUT_4</name></connection>
<connection>
<GID>688</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-29.5,615,-29.5</points>
<connection>
<GID>686</GID>
<name>OUT_3</name></connection>
<connection>
<GID>688</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-30.5,615,-30.5</points>
<connection>
<GID>686</GID>
<name>OUT_2</name></connection>
<connection>
<GID>688</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-31.5,615,-31.5</points>
<connection>
<GID>686</GID>
<name>OUT_1</name></connection>
<connection>
<GID>688</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>606,-32.5,615,-32.5</points>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection>
<connection>
<GID>688</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-25.5,629,-25.5</points>
<connection>
<GID>688</GID>
<name>OUT_7</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-26.5,629,-26.5</points>
<connection>
<GID>688</GID>
<name>OUT_6</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-27.5,629,-27.5</points>
<connection>
<GID>688</GID>
<name>OUT_5</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-28.5,629,-28.5</points>
<connection>
<GID>688</GID>
<name>OUT_4</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-29.5,629,-29.5</points>
<connection>
<GID>688</GID>
<name>OUT_3</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-30.5,629,-30.5</points>
<connection>
<GID>688</GID>
<name>OUT_2</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,-23.5,618,-13</points>
<connection>
<GID>688</GID>
<name>load</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>615,-13,618,-13</points>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection>
<intersection>618 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>602,-23.5,602,-10.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<connection>
<GID>686</GID>
<name>count_enable</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>602,-22.5,603,-22.5</points>
<intersection>602 0</intersection>
<intersection>603 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>603,-23.5,603,-22.5</points>
<connection>
<GID>686</GID>
<name>count_up</name></connection>
<intersection>-22.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>656,-62,656,-60.5</points>
<connection>
<GID>690</GID>
<name>load</name></connection>
<intersection>-60.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>655.5,-60.5,656,-60.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>656 3</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-31.5,629,-31.5</points>
<connection>
<GID>688</GID>
<name>OUT_1</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-32.5,629,-32.5</points>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-64,670.5,-64</points>
<connection>
<GID>690</GID>
<name>OUT_7</name></connection>
<connection>
<GID>692</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-65,670.5,-65</points>
<connection>
<GID>690</GID>
<name>OUT_6</name></connection>
<connection>
<GID>692</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-66,670.5,-66</points>
<connection>
<GID>690</GID>
<name>OUT_5</name></connection>
<connection>
<GID>692</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-67,670.5,-67</points>
<connection>
<GID>690</GID>
<name>OUT_4</name></connection>
<connection>
<GID>692</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-68,670.5,-68</points>
<connection>
<GID>690</GID>
<name>OUT_3</name></connection>
<connection>
<GID>692</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-69,670.5,-69</points>
<connection>
<GID>690</GID>
<name>OUT_2</name></connection>
<connection>
<GID>692</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-70,670.5,-70</points>
<connection>
<GID>690</GID>
<name>OUT_1</name></connection>
<connection>
<GID>692</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-71,670.5,-71</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<connection>
<GID>692</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673.5,-62,673.5,-60.5</points>
<connection>
<GID>692</GID>
<name>load</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>673,-60.5,673.5,-60.5</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<intersection>673.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>678.5,-71,682,-71</points>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection>
<connection>
<GID>708</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>678.5,-70,682,-70</points>
<connection>
<GID>692</GID>
<name>OUT_1</name></connection>
<connection>
<GID>708</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,-59,618,-34.5</points>
<connection>
<GID>688</GID>
<name>clock</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-59,666,-59</points>
<intersection>585.5 10</intersection>
<intersection>588 6</intersection>
<intersection>618 0</intersection>
<intersection>651.5 5</intersection>
<intersection>666 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>666,-73,666,-59</points>
<intersection>-73 11</intersection>
<intersection>-59 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>651.5,-73.5,651.5,-59</points>
<intersection>-73.5 8</intersection>
<intersection>-59 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>588,-59,588,-41.5</points>
<intersection>-59 1</intersection>
<intersection>-41.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>588,-41.5,594,-41.5</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>588 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>651.5,-73.5,656,-73.5</points>
<intersection>651.5 5</intersection>
<intersection>656 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>656,-73.5,656,-73</points>
<connection>
<GID>690</GID>
<name>clock</name></connection>
<intersection>-73.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>585.5,-60,585.5,-59</points>
<connection>
<GID>719</GID>
<name>OUT</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>666,-73,673.5,-73</points>
<connection>
<GID>692</GID>
<name>clock</name></connection>
<intersection>666 4</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-58.5,603,-34.5</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<connection>
<GID>686</GID>
<name>clear</name></connection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>603,-58.5,665.5,-58.5</points>
<intersection>603 0</intersection>
<intersection>620 3</intersection>
<intersection>651 7</intersection>
<intersection>665.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>620,-58.5,620,-34.5</points>
<connection>
<GID>688</GID>
<name>clear</name></connection>
<intersection>-58.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>665.5,-73.5,665.5,-58.5</points>
<intersection>-73.5 10</intersection>
<intersection>-58.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>651,-74,651,-58.5</points>
<intersection>-74 8</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>651,-74,658,-74</points>
<intersection>651 7</intersection>
<intersection>658 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>658,-74,658,-73</points>
<connection>
<GID>690</GID>
<name>clear</name></connection>
<intersection>-74 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>665.5,-73.5,675.5,-73.5</points>
<intersection>665.5 6</intersection>
<intersection>675.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>675.5,-73.5,675.5,-73</points>
<connection>
<GID>692</GID>
<name>clear</name></connection>
<intersection>-73.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,-26.5,642,-26.5</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>640 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>640,-41.5,640,-26.5</points>
<intersection>-41.5 4</intersection>
<intersection>-28.5 7</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>625.5,-41.5,640,-41.5</points>
<intersection>625.5 8</intersection>
<intersection>640 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>639,-28.5,640,-28.5</points>
<connection>
<GID>691</GID>
<name>write_enable</name></connection>
<intersection>640 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>625.5,-62.5,625.5,-41.5</points>
<connection>
<GID>714</GID>
<name>ENABLE_0</name></connection>
<intersection>-41.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>639,-29.5,642,-29.5</points>
<connection>
<GID>691</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>710</GID>
<name>OUT_0</name></connection>
<intersection>642 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>642,-41.5,642,-29.5</points>
<intersection>-41.5 6</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>642,-41.5,647.5,-41.5</points>
<intersection>642 5</intersection>
<intersection>647.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>647.5,-62.5,647.5,-41.5</points>
<connection>
<GID>713</GID>
<name>ENABLE_0</name></connection>
<intersection>-41.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-70,645.5,-70</points>
<connection>
<GID>714</GID>
<name>OUT_1</name></connection>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>636.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>636.5,-70,636.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_1</name></connection>
<intersection>-70 1</intersection></vsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-69,645.5,-69</points>
<connection>
<GID>714</GID>
<name>OUT_2</name></connection>
<connection>
<GID>713</GID>
<name>IN_2</name></connection>
<intersection>635.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>635.5,-69,635.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_2</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-68,645.5,-68</points>
<connection>
<GID>714</GID>
<name>OUT_3</name></connection>
<connection>
<GID>713</GID>
<name>IN_3</name></connection>
<intersection>634.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>634.5,-68,634.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_3</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-67,645.5,-67</points>
<connection>
<GID>714</GID>
<name>OUT_4</name></connection>
<connection>
<GID>713</GID>
<name>IN_4</name></connection>
<intersection>633.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>633.5,-67,633.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_4</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-66,645.5,-66</points>
<connection>
<GID>714</GID>
<name>OUT_5</name></connection>
<connection>
<GID>713</GID>
<name>IN_5</name></connection>
<intersection>632.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>632.5,-66,632.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_5</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-65,645.5,-65</points>
<connection>
<GID>714</GID>
<name>OUT_6</name></connection>
<connection>
<GID>713</GID>
<name>IN_6</name></connection>
<intersection>631.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>631.5,-65,631.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_6</name></connection>
<intersection>-65 1</intersection></vsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-64,645.5,-64</points>
<connection>
<GID>714</GID>
<name>OUT_7</name></connection>
<connection>
<GID>713</GID>
<name>IN_7</name></connection>
<intersection>630.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>630.5,-64,630.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_7</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-66,653,-66</points>
<connection>
<GID>713</GID>
<name>OUT_5</name></connection>
<connection>
<GID>690</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-71,653,-71</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<connection>
<GID>690</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-70,653,-70</points>
<connection>
<GID>713</GID>
<name>OUT_1</name></connection>
<connection>
<GID>690</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-69,653,-69</points>
<connection>
<GID>713</GID>
<name>OUT_2</name></connection>
<connection>
<GID>690</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-68,653,-68</points>
<connection>
<GID>713</GID>
<name>OUT_3</name></connection>
<connection>
<GID>690</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-67,653,-67</points>
<connection>
<GID>713</GID>
<name>OUT_4</name></connection>
<connection>
<GID>690</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-64,653,-64</points>
<connection>
<GID>713</GID>
<name>OUT_7</name></connection>
<connection>
<GID>690</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-65,653,-65</points>
<connection>
<GID>713</GID>
<name>OUT_6</name></connection>
<connection>
<GID>690</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-71,645.5,-71</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>637.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>637.5,-71,637.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>692,-68,694,-68</points>
<connection>
<GID>708</GID>
<name>ENABLE_0</name></connection>
<intersection>694 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>694,-68,694,-47</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>575,-61,579.5,-61</points>
<connection>
<GID>695</GID>
<name>CLK</name></connection>
<connection>
<GID>719</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579.5,-59,579.5,-57</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>579,-57,579.5,-57</points>
<connection>
<GID>720</GID>
<name>OUT_0</name></connection>
<intersection>579.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601,-42.5,601,-34.5</points>
<connection>
<GID>686</GID>
<name>clock</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>600,-42.5,601,-42.5</points>
<connection>
<GID>718</GID>
<name>OUT</name></connection>
<intersection>601 0</intersection></hsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>570,-43.5,594,-43.5</points>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection>
<connection>
<GID>718</GID>
<name>IN_1</name></connection>
<intersection>573 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>573,-43.5,573,-41</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601,-23.5,601,-15.5</points>
<connection>
<GID>686</GID>
<name>load</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>573,-35,573,-15.5</points>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>573,-15.5,601,-15.5</points>
<intersection>573 1</intersection>
<intersection>601 0</intersection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>626,-84,626,-84</points>
<connection>
<GID>770</GID>
<name>ENABLE</name></connection>
<connection>
<GID>771</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>605,-78.5,661,-78.5</points>
<intersection>605 8</intersection>
<intersection>661 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>661,-130,661,-78.5</points>
<intersection>-130 18</intersection>
<intersection>-125 19</intersection>
<intersection>-120 20</intersection>
<intersection>-115 21</intersection>
<intersection>-110 22</intersection>
<intersection>-105 23</intersection>
<intersection>-100 24</intersection>
<intersection>-95 25</intersection>
<intersection>-78.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>605,-87,605,-78.5</points>
<intersection>-87 10</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>605,-87,626,-87</points>
<connection>
<GID>772</GID>
<name>OUT_0</name></connection>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>605 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>661,-130,680.5,-130</points>
<connection>
<GID>798</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>661,-125,680.5,-125</points>
<connection>
<GID>797</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>661,-120,680.5,-120</points>
<connection>
<GID>796</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>661,-115,680.5,-115</points>
<connection>
<GID>795</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>661,-110,680.5,-110</points>
<connection>
<GID>794</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>661,-105,680.5,-105</points>
<connection>
<GID>793</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>661,-100,680.5,-100</points>
<connection>
<GID>792</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>661,-95,680.5,-95</points>
<connection>
<GID>791</GID>
<name>SEL_0</name></connection>
<intersection>661 7</intersection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>633,-116,633,-87</points>
<intersection>-116 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>632,-87,633,-87</points>
<connection>
<GID>770</GID>
<name>OUT_0</name></connection>
<intersection>633 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>633,-116,637.5,-116</points>
<connection>
<GID>723</GID>
<name>ENABLE_0</name></connection>
<intersection>633 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>637.5,-93,637.5,-86</points>
<connection>
<GID>722</GID>
<name>ENABLE_0</name></connection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>632,-86,637.5,-86</points>
<connection>
<GID>770</GID>
<name>OUT_1</name></connection>
<intersection>637.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>654,-129,654,-129</points>
<connection>
<GID>775</GID>
<name>carry_out</name></connection>
<connection>
<GID>776</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641,-132.5,641,-116</points>
<intersection>-132.5 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641,-116,651,-116</points>
<connection>
<GID>775</GID>
<name>IN_B_0</name></connection>
<intersection>641 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-132.5,641,-132.5</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>641 0</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641.5,-130.5,641.5,-117</points>
<intersection>-130.5 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641.5,-117,651,-117</points>
<connection>
<GID>775</GID>
<name>IN_B_1</name></connection>
<intersection>641.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-130.5,641.5,-130.5</points>
<connection>
<GID>723</GID>
<name>OUT_2</name></connection>
<intersection>641.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642,-128.5,642,-118</points>
<intersection>-128.5 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642,-118,651,-118</points>
<connection>
<GID>775</GID>
<name>IN_B_2</name></connection>
<intersection>642 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-128.5,642,-128.5</points>
<connection>
<GID>723</GID>
<name>OUT_4</name></connection>
<intersection>642 0</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642.5,-126.5,642.5,-119</points>
<intersection>-126.5 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642.5,-119,651,-119</points>
<connection>
<GID>775</GID>
<name>IN_B_3</name></connection>
<intersection>642.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-126.5,642.5,-126.5</points>
<connection>
<GID>723</GID>
<name>OUT_6</name></connection>
<intersection>642.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644.5,-132,644.5,-124.5</points>
<intersection>-132 1</intersection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644.5,-132,651,-132</points>
<connection>
<GID>776</GID>
<name>IN_B_0</name></connection>
<intersection>644.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-124.5,644.5,-124.5</points>
<connection>
<GID>723</GID>
<name>OUT_8</name></connection>
<intersection>644.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-133,644,-122.5</points>
<intersection>-133 1</intersection>
<intersection>-122.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-133,651,-133</points>
<connection>
<GID>776</GID>
<name>IN_B_1</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-122.5,644,-122.5</points>
<connection>
<GID>723</GID>
<name>OUT_10</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643.5,-134,643.5,-120.5</points>
<intersection>-134 1</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643.5,-134,651,-134</points>
<connection>
<GID>776</GID>
<name>IN_B_2</name></connection>
<intersection>643.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-120.5,643.5,-120.5</points>
<connection>
<GID>723</GID>
<name>OUT_12</name></connection>
<intersection>643.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643,-135,643,-118.5</points>
<intersection>-135 1</intersection>
<intersection>-118.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643,-135,651,-135</points>
<connection>
<GID>776</GID>
<name>IN_B_3</name></connection>
<intersection>643 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-118.5,643,-118.5</points>
<connection>
<GID>723</GID>
<name>OUT_14</name></connection>
<intersection>643 0</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,-131.5,645,-123</points>
<intersection>-131.5 2</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645,-123,651,-123</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>645 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-131.5,645,-131.5</points>
<connection>
<GID>723</GID>
<name>OUT_1</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,-129.5,645,-124</points>
<intersection>-129.5 2</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645,-124,651,-124</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>645 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-129.5,645,-129.5</points>
<connection>
<GID>723</GID>
<name>OUT_3</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,-127.5,645,-125</points>
<intersection>-127.5 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645,-125,651,-125</points>
<connection>
<GID>775</GID>
<name>IN_2</name></connection>
<intersection>645 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-127.5,645,-127.5</points>
<connection>
<GID>723</GID>
<name>OUT_5</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,-126,645,-125.5</points>
<intersection>-126 1</intersection>
<intersection>-125.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645,-126,651,-126</points>
<connection>
<GID>775</GID>
<name>IN_3</name></connection>
<intersection>645 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-125.5,645,-125.5</points>
<connection>
<GID>723</GID>
<name>OUT_7</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>647,-139,647,-123.5</points>
<intersection>-139 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>647,-139,651,-139</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>647 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-123.5,647,-123.5</points>
<connection>
<GID>723</GID>
<name>OUT_9</name></connection>
<intersection>647 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646.5,-140,646.5,-121.5</points>
<intersection>-140 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646.5,-140,651,-140</points>
<connection>
<GID>776</GID>
<name>IN_1</name></connection>
<intersection>646.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-121.5,646.5,-121.5</points>
<connection>
<GID>723</GID>
<name>OUT_11</name></connection>
<intersection>646.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646,-141,646,-119.5</points>
<intersection>-141 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,-141,651,-141</points>
<connection>
<GID>776</GID>
<name>IN_2</name></connection>
<intersection>646 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-119.5,646,-119.5</points>
<connection>
<GID>723</GID>
<name>OUT_13</name></connection>
<intersection>646 0</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645.5,-142,645.5,-117.5</points>
<intersection>-142 1</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645.5,-142,651,-142</points>
<connection>
<GID>776</GID>
<name>IN_3</name></connection>
<intersection>645.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-117.5,645.5,-117.5</points>
<connection>
<GID>723</GID>
<name>OUT_15</name></connection>
<intersection>645.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>647,-111.5,647.5,-111.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>647 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>647,-111.5,647,-109.5</points>
<intersection>-111.5 1</intersection>
<intersection>-109.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>639.5,-109.5,647,-109.5</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>647 3</intersection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>639.5,-108.5,646.5,-108.5</points>
<connection>
<GID>722</GID>
<name>OUT_1</name></connection>
<intersection>646.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>646.5,-109.5,646.5,-108.5</points>
<intersection>-109.5 5</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>646.5,-109.5,647.5,-109.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>646.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646,-108,646,-107.5</points>
<intersection>-108 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,-108,652.5,-108</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>646 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-107.5,646,-107.5</points>
<connection>
<GID>722</GID>
<name>OUT_2</name></connection>
<intersection>646 0</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>639.5,-106.5,652.5,-106.5</points>
<connection>
<GID>722</GID>
<name>OUT_3</name></connection>
<intersection>652.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>652.5,-106.5,652.5,-106</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>-106.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>639.5,-105.5,647.5,-105.5</points>
<connection>
<GID>722</GID>
<name>OUT_4</name></connection>
<intersection>647.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>647.5,-105.5,647.5,-104.5</points>
<connection>
<GID>785</GID>
<name>IN_1</name></connection>
<intersection>-105.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644.5,-104.5,644.5,-102.5</points>
<intersection>-104.5 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644.5,-102.5,647.5,-102.5</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>644.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-104.5,644.5,-104.5</points>
<connection>
<GID>722</GID>
<name>OUT_5</name></connection>
<intersection>644.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-103.5,644,-101</points>
<intersection>-103.5 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-101,652.5,-101</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-103.5,644,-103.5</points>
<connection>
<GID>722</GID>
<name>OUT_6</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643.5,-102.5,643.5,-99</points>
<intersection>-102.5 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643.5,-99,652.5,-99</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>643.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-102.5,643.5,-102.5</points>
<connection>
<GID>722</GID>
<name>OUT_7</name></connection>
<intersection>643.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643,-101.5,643,-97.5</points>
<intersection>-101.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643,-97.5,647.5,-97.5</points>
<connection>
<GID>787</GID>
<name>IN_1</name></connection>
<intersection>643 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-101.5,643,-101.5</points>
<connection>
<GID>722</GID>
<name>OUT_8</name></connection>
<intersection>643 0</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642.5,-100.5,642.5,-95.5</points>
<intersection>-100.5 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642.5,-95.5,647.5,-95.5</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>642.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-100.5,642.5,-100.5</points>
<connection>
<GID>722</GID>
<name>OUT_9</name></connection>
<intersection>642.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642,-99.5,642,-94</points>
<intersection>-99.5 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642,-94,652.5,-94</points>
<connection>
<GID>788</GID>
<name>IN_1</name></connection>
<intersection>642 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-99.5,642,-99.5</points>
<connection>
<GID>722</GID>
<name>OUT_10</name></connection>
<intersection>642 0</intersection></hsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641.5,-98.5,641.5,-92</points>
<intersection>-98.5 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641.5,-92,652.5,-92</points>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>641.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-98.5,641.5,-98.5</points>
<connection>
<GID>722</GID>
<name>OUT_11</name></connection>
<intersection>641.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641,-97.5,641,-90.5</points>
<intersection>-97.5 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641,-90.5,647.5,-90.5</points>
<connection>
<GID>789</GID>
<name>IN_1</name></connection>
<intersection>641 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-97.5,641,-97.5</points>
<connection>
<GID>722</GID>
<name>OUT_12</name></connection>
<intersection>641 0</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640.5,-96.5,640.5,-88.5</points>
<intersection>-96.5 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640.5,-88.5,647.5,-88.5</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>640.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-96.5,640.5,-96.5</points>
<connection>
<GID>722</GID>
<name>OUT_13</name></connection>
<intersection>640.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,-95.5,640,-87</points>
<intersection>-95.5 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,-87,652.5,-87</points>
<connection>
<GID>790</GID>
<name>IN_1</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,-95.5,640,-95.5</points>
<connection>
<GID>722</GID>
<name>OUT_14</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-94.5,639.5,-85</points>
<connection>
<GID>722</GID>
<name>OUT_15</name></connection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-85,652.5,-85</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-133.5,668.5,-119.5</points>
<intersection>-133.5 1</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-133.5,678.5,-133.5</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-119.5,668.5,-119.5</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-128.5,668.5,-120.5</points>
<intersection>-128.5 1</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-128.5,678.5,-128.5</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-120.5,668.5,-120.5</points>
<connection>
<GID>775</GID>
<name>OUT_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-123.5,668.5,-121.5</points>
<intersection>-123.5 1</intersection>
<intersection>-121.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-123.5,678.5,-123.5</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-121.5,668.5,-121.5</points>
<connection>
<GID>775</GID>
<name>OUT_2</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-122.5,668.5,-118.5</points>
<intersection>-122.5 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-118.5,678.5,-118.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-122.5,668.5,-122.5</points>
<connection>
<GID>775</GID>
<name>OUT_3</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-135.5,668.5,-113.5</points>
<intersection>-135.5 2</intersection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-113.5,678.5,-113.5</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-135.5,668.5,-135.5</points>
<connection>
<GID>776</GID>
<name>OUT_0</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-136.5,668.5,-108.5</points>
<intersection>-136.5 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-108.5,678.5,-108.5</points>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-136.5,668.5,-136.5</points>
<connection>
<GID>776</GID>
<name>OUT_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-137.5,668.5,-103.5</points>
<intersection>-137.5 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-103.5,678.5,-103.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-137.5,668.5,-137.5</points>
<connection>
<GID>776</GID>
<name>OUT_2</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-138.5,668.5,-98.5</points>
<intersection>-138.5 2</intersection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>668.5,-98.5,678.5,-98.5</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>659,-138.5,668.5,-138.5</points>
<connection>
<GID>776</GID>
<name>OUT_3</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,-131.5,666,-110.5</points>
<intersection>-131.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>666,-131.5,678.5,-131.5</points>
<connection>
<GID>798</GID>
<name>IN_1</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>653.5,-110.5,666,-110.5</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-126.5,668.5,-107</points>
<intersection>-126.5 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>658.5,-107,668.5,-107</points>
<connection>
<GID>784</GID>
<name>OUT</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>668.5,-126.5,678.5,-126.5</points>
<connection>
<GID>797</GID>
<name>IN_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,-121.5,666,-103.5</points>
<intersection>-121.5 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-103.5,666,-103.5</points>
<connection>
<GID>785</GID>
<name>OUT</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>666,-121.5,678.5,-121.5</points>
<connection>
<GID>796</GID>
<name>IN_1</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-116.5,668.5,-100</points>
<intersection>-116.5 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>658.5,-100,668.5,-100</points>
<connection>
<GID>786</GID>
<name>OUT</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>668.5,-116.5,678.5,-116.5</points>
<connection>
<GID>795</GID>
<name>IN_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,-111.5,666,-96.5</points>
<intersection>-111.5 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-96.5,666,-96.5</points>
<connection>
<GID>787</GID>
<name>OUT</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>666,-111.5,678.5,-111.5</points>
<connection>
<GID>794</GID>
<name>IN_1</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-106.5,668.5,-93</points>
<intersection>-106.5 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>658.5,-93,668.5,-93</points>
<connection>
<GID>788</GID>
<name>OUT</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>668.5,-106.5,678.5,-106.5</points>
<connection>
<GID>793</GID>
<name>IN_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,-101.5,666,-89.5</points>
<intersection>-101.5 2</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-89.5,666,-89.5</points>
<connection>
<GID>789</GID>
<name>OUT</name></connection>
<intersection>666 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>666,-101.5,678.5,-101.5</points>
<connection>
<GID>792</GID>
<name>IN_1</name></connection>
<intersection>666 0</intersection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,-96.5,668.5,-86</points>
<intersection>-96.5 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>658.5,-86,668.5,-86</points>
<connection>
<GID>790</GID>
<name>OUT</name></connection>
<intersection>668.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>668.5,-96.5,678.5,-96.5</points>
<connection>
<GID>791</GID>
<name>IN_1</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-132.5,690,-117.5</points>
<intersection>-132.5 2</intersection>
<intersection>-117.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-117.5,698,-117.5</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>690 0</intersection>
<intersection>691 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-132.5,690,-132.5</points>
<connection>
<GID>798</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>691,-123,691,-117.5</points>
<intersection>-123 8</intersection>
<intersection>-117.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>691,-123,712,-123</points>
<intersection>691 7</intersection>
<intersection>712 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>712,-123.5,712,-123</points>
<connection>
<GID>809</GID>
<name>N_in2</name></connection>
<intersection>-123 8</intersection></vsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-127.5,690,-116.5</points>
<intersection>-127.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-116.5,698,-116.5</points>
<connection>
<GID>799</GID>
<name>IN_1</name></connection>
<intersection>690 0</intersection>
<intersection>691.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-127.5,690,-127.5</points>
<connection>
<GID>797</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>691.5,-122.5,691.5,-116.5</points>
<intersection>-122.5 8</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>691.5,-122.5,709.5,-122.5</points>
<intersection>691.5 7</intersection>
<intersection>709.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>709.5,-123.5,709.5,-122.5</points>
<connection>
<GID>808</GID>
<name>N_in2</name></connection>
<intersection>-122.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-122.5,690,-115.5</points>
<intersection>-122.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-115.5,698,-115.5</points>
<connection>
<GID>799</GID>
<name>IN_2</name></connection>
<intersection>690 0</intersection>
<intersection>692 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-122.5,690,-122.5</points>
<connection>
<GID>796</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>692,-122,692,-115.5</points>
<intersection>-122 8</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>692,-122,707,-122</points>
<intersection>692 7</intersection>
<intersection>707 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>707,-123.5,707,-122</points>
<connection>
<GID>807</GID>
<name>N_in2</name></connection>
<intersection>-122 8</intersection></vsegment></shape></wire>
<wire>
<ID>1140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-117.5,690,-114.5</points>
<intersection>-117.5 2</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-114.5,698,-114.5</points>
<connection>
<GID>799</GID>
<name>IN_3</name></connection>
<intersection>690 0</intersection>
<intersection>692.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-117.5,690,-117.5</points>
<connection>
<GID>795</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>692.5,-121.5,692.5,-114.5</points>
<intersection>-121.5 9</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>692.5,-121.5,704.5,-121.5</points>
<intersection>692.5 8</intersection>
<intersection>704.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>704.5,-123.5,704.5,-121.5</points>
<connection>
<GID>806</GID>
<name>N_in2</name></connection>
<intersection>-121.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>1141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-113.5,690,-112.5</points>
<intersection>-113.5 1</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-113.5,698,-113.5</points>
<connection>
<GID>799</GID>
<name>IN_4</name></connection>
<intersection>690 0</intersection>
<intersection>693 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-112.5,690,-112.5</points>
<connection>
<GID>794</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>693,-121,693,-113.5</points>
<intersection>-121 9</intersection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>693,-121,702,-121</points>
<intersection>693 8</intersection>
<intersection>702 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>702,-123.5,702,-121</points>
<connection>
<GID>805</GID>
<name>N_in2</name></connection>
<intersection>-121 9</intersection></vsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-112.5,690,-107.5</points>
<intersection>-112.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-112.5,698,-112.5</points>
<connection>
<GID>799</GID>
<name>IN_5</name></connection>
<intersection>690 0</intersection>
<intersection>693.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-107.5,690,-107.5</points>
<connection>
<GID>793</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>693.5,-120.5,693.5,-112.5</points>
<intersection>-120.5 8</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>693.5,-120.5,699.5,-120.5</points>
<intersection>693.5 7</intersection>
<intersection>699.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>699.5,-123.5,699.5,-120.5</points>
<connection>
<GID>804</GID>
<name>N_in2</name></connection>
<intersection>-120.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-111.5,690,-102.5</points>
<intersection>-111.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>690,-111.5,698,-111.5</points>
<connection>
<GID>799</GID>
<name>IN_6</name></connection>
<intersection>690 0</intersection>
<intersection>694 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>682.5,-102.5,690,-102.5</points>
<connection>
<GID>792</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>694,-120,694,-111.5</points>
<intersection>-120 8</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>694,-120,697,-120</points>
<intersection>694 7</intersection>
<intersection>697 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>697,-123.5,697,-120</points>
<connection>
<GID>803</GID>
<name>N_in2</name></connection>
<intersection>-120 8</intersection></vsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597,-152,597,-150</points>
<intersection>-152 2</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,-150,624.5,-150</points>
<connection>
<GID>129</GID>
<name>IN_15</name></connection>
<intersection>597 0</intersection>
<intersection>599.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-152,597,-152</points>
<connection>
<GID>132</GID>
<name>OUT_7</name></connection>
<intersection>597 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>599.5,-173,599.5,-150</points>
<intersection>-173 4</intersection>
<intersection>-150 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>599.5,-173,624.5,-173</points>
<connection>
<GID>130</GID>
<name>IN_15</name></connection>
<intersection>599.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-110.5,690,-97.5</points>
<intersection>-110.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>682.5,-97.5,690,-97.5</points>
<connection>
<GID>791</GID>
<name>OUT</name></connection>
<intersection>690 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>690,-110.5,698,-110.5</points>
<connection>
<GID>799</GID>
<name>IN_7</name></connection>
<intersection>690 0</intersection>
<intersection>694.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>694.5,-123.5,694.5,-110.5</points>
<connection>
<GID>802</GID>
<name>N_in2</name></connection>
<intersection>-110.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597.5,-153,597.5,-152</points>
<intersection>-153 2</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597.5,-152,624.5,-152</points>
<connection>
<GID>129</GID>
<name>IN_13</name></connection>
<intersection>597.5 0</intersection>
<intersection>600.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-153,597.5,-153</points>
<connection>
<GID>132</GID>
<name>OUT_6</name></connection>
<intersection>597.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>600.5,-175,600.5,-152</points>
<intersection>-175 4</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>600.5,-175,624.5,-175</points>
<connection>
<GID>130</GID>
<name>IN_13</name></connection>
<intersection>600.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-85,503.5,-85</points>
<connection>
<GID>687</GID>
<name>OUT_7</name></connection>
<intersection>503.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>503.5,-85,503.5,-75</points>
<intersection>-85 1</intersection>
<intersection>-75 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503.5,-75,534,-75</points>
<connection>
<GID>727</GID>
<name>IN_3</name></connection>
<connection>
<GID>744</GID>
<name>IN_3</name></connection>
<intersection>503.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>588.5,-154,624.5,-154</points>
<connection>
<GID>132</GID>
<name>OUT_5</name></connection>
<connection>
<GID>129</GID>
<name>IN_11</name></connection>
<intersection>601.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>601.5,-177,601.5,-154</points>
<intersection>-177 3</intersection>
<intersection>-154 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>601.5,-177,624.5,-177</points>
<connection>
<GID>130</GID>
<name>IN_11</name></connection>
<intersection>601.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-86,534,-86</points>
<connection>
<GID>687</GID>
<name>OUT_6</name></connection>
<connection>
<GID>728</GID>
<name>IN_3</name></connection>
<connection>
<GID>745</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597,-156,597,-155</points>
<intersection>-156 1</intersection>
<intersection>-155 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,-156,624.5,-156</points>
<connection>
<GID>129</GID>
<name>IN_9</name></connection>
<intersection>597 0</intersection>
<intersection>602.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-155,597,-155</points>
<connection>
<GID>132</GID>
<name>OUT_4</name></connection>
<intersection>597 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>602.5,-179,602.5,-156</points>
<intersection>-179 4</intersection>
<intersection>-156 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>602.5,-179,624.5,-179</points>
<connection>
<GID>130</GID>
<name>IN_9</name></connection>
<intersection>602.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504.5,-97,504.5,-87</points>
<intersection>-97 1</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504.5,-97,534,-97</points>
<connection>
<GID>729</GID>
<name>IN_3</name></connection>
<connection>
<GID>746</GID>
<name>IN_3</name></connection>
<intersection>504.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-87,504.5,-87</points>
<connection>
<GID>687</GID>
<name>OUT_5</name></connection>
<intersection>504.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,-158,596.5,-156</points>
<intersection>-158 1</intersection>
<intersection>-156 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596.5,-158,624.5,-158</points>
<connection>
<GID>129</GID>
<name>IN_7</name></connection>
<intersection>596.5 0</intersection>
<intersection>603.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-156,596.5,-156</points>
<connection>
<GID>132</GID>
<name>OUT_3</name></connection>
<intersection>596.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>603.5,-181,603.5,-158</points>
<intersection>-181 4</intersection>
<intersection>-158 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>603.5,-181,624.5,-181</points>
<connection>
<GID>130</GID>
<name>IN_7</name></connection>
<intersection>603.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505,-106.5,505,-88</points>
<intersection>-106.5 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505,-106.5,534,-106.5</points>
<connection>
<GID>747</GID>
<name>IN_3</name></connection>
<connection>
<GID>730</GID>
<name>IN_3</name></connection>
<intersection>505 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-88,505,-88</points>
<connection>
<GID>687</GID>
<name>OUT_4</name></connection>
<intersection>505 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596,-160,596,-157</points>
<intersection>-160 1</intersection>
<intersection>-157 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596,-160,624.5,-160</points>
<connection>
<GID>129</GID>
<name>IN_5</name></connection>
<intersection>596 0</intersection>
<intersection>604.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-157,596,-157</points>
<connection>
<GID>132</GID>
<name>OUT_2</name></connection>
<intersection>596 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>604.5,-183,604.5,-160</points>
<intersection>-183 4</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>604.5,-183,624.5,-183</points>
<connection>
<GID>130</GID>
<name>IN_5</name></connection>
<intersection>604.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,-117.5,505.5,-89</points>
<intersection>-117.5 1</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505.5,-117.5,534,-117.5</points>
<connection>
<GID>731</GID>
<name>IN_3</name></connection>
<connection>
<GID>748</GID>
<name>IN_3</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-89,505.5,-89</points>
<connection>
<GID>687</GID>
<name>OUT_3</name></connection>
<intersection>505.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>595.5,-162,595.5,-158</points>
<intersection>-162 1</intersection>
<intersection>-158 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595.5,-162,624.5,-162</points>
<connection>
<GID>129</GID>
<name>IN_3</name></connection>
<intersection>595.5 0</intersection>
<intersection>605.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-158,595.5,-158</points>
<connection>
<GID>132</GID>
<name>OUT_1</name></connection>
<intersection>595.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>605.5,-185,605.5,-162</points>
<intersection>-185 4</intersection>
<intersection>-162 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>605.5,-185,624.5,-185</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>605.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506,-128.5,506,-90</points>
<intersection>-128.5 1</intersection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>506,-128.5,534,-128.5</points>
<connection>
<GID>732</GID>
<name>IN_3</name></connection>
<connection>
<GID>749</GID>
<name>IN_3</name></connection>
<intersection>506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-90,506,-90</points>
<connection>
<GID>687</GID>
<name>OUT_2</name></connection>
<intersection>506 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>595,-164,595,-159</points>
<intersection>-164 1</intersection>
<intersection>-159 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595,-164,624.5,-164</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>595 0</intersection>
<intersection>606.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-159,595,-159</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>595 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>606.5,-187,606.5,-164</points>
<intersection>-187 4</intersection>
<intersection>-164 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>606.5,-187,624.5,-187</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>606.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-139,508,-91</points>
<intersection>-139 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-139,534,-139</points>
<connection>
<GID>733</GID>
<name>IN_3</name></connection>
<connection>
<GID>750</GID>
<name>IN_3</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-91,508,-91</points>
<connection>
<GID>687</GID>
<name>OUT_1</name></connection>
<intersection>508 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-183.5,589.5,-174</points>
<intersection>-183.5 2</intersection>
<intersection>-174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,-174,624.5,-174</points>
<connection>
<GID>130</GID>
<name>IN_14</name></connection>
<intersection>589.5 0</intersection>
<intersection>600 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-183.5,589.5,-183.5</points>
<connection>
<GID>134</GID>
<name>OUT_7</name></connection>
<intersection>589.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>600,-174,600,-151</points>
<intersection>-174 1</intersection>
<intersection>-151 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>600,-151,624.5,-151</points>
<connection>
<GID>129</GID>
<name>IN_14</name></connection>
<intersection>600 3</intersection></hsegment></shape></wire>
<wire>
<ID>1152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>507,-150,507,-92</points>
<intersection>-150 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,-92,507,-92</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>507 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>507,-150,534,-150</points>
<connection>
<GID>734</GID>
<name>IN_3</name></connection>
<connection>
<GID>751</GID>
<name>IN_3</name></connection>
<intersection>507 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,-184.5,590,-176</points>
<intersection>-184.5 2</intersection>
<intersection>-176 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,-176,624.5,-176</points>
<connection>
<GID>130</GID>
<name>IN_12</name></connection>
<intersection>590 0</intersection>
<intersection>601 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-184.5,590,-184.5</points>
<connection>
<GID>134</GID>
<name>OUT_6</name></connection>
<intersection>590 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>601,-176,601,-153</points>
<intersection>-176 1</intersection>
<intersection>-153 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>601,-153,624.5,-153</points>
<connection>
<GID>129</GID>
<name>IN_12</name></connection>
<intersection>601 3</intersection></hsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508,-98,508,-77</points>
<intersection>-98 2</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,-77,534,-77</points>
<connection>
<GID>744</GID>
<name>IN_2</name></connection>
<connection>
<GID>727</GID>
<name>IN_2</name></connection>
<intersection>508 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-98,508,-98</points>
<connection>
<GID>689</GID>
<name>OUT_7</name></connection>
<intersection>508 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,-185.5,590.5,-178</points>
<intersection>-185.5 2</intersection>
<intersection>-178 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,-178,624.5,-178</points>
<connection>
<GID>130</GID>
<name>IN_10</name></connection>
<intersection>590.5 0</intersection>
<intersection>602 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-185.5,590.5,-185.5</points>
<connection>
<GID>134</GID>
<name>OUT_5</name></connection>
<intersection>590.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>602,-178,602,-155</points>
<intersection>-178 1</intersection>
<intersection>-155 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>602,-155,624.5,-155</points>
<connection>
<GID>129</GID>
<name>IN_10</name></connection>
<intersection>602 3</intersection></hsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>508.5,-99,508.5,-88</points>
<intersection>-99 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508.5,-88,534,-88</points>
<connection>
<GID>728</GID>
<name>IN_2</name></connection>
<connection>
<GID>745</GID>
<name>IN_2</name></connection>
<intersection>508.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-99,508.5,-99</points>
<connection>
<GID>689</GID>
<name>OUT_6</name></connection>
<intersection>508.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591,-186.5,591,-180</points>
<intersection>-186.5 2</intersection>
<intersection>-180 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591,-180,624.5,-180</points>
<connection>
<GID>130</GID>
<name>IN_8</name></connection>
<intersection>591 0</intersection>
<intersection>603 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-186.5,591,-186.5</points>
<connection>
<GID>134</GID>
<name>OUT_4</name></connection>
<intersection>591 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>603,-180,603,-157</points>
<intersection>-180 1</intersection>
<intersection>-157 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>603,-157,624.5,-157</points>
<connection>
<GID>129</GID>
<name>IN_8</name></connection>
<intersection>603 3</intersection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-100,509,-100</points>
<connection>
<GID>689</GID>
<name>OUT_5</name></connection>
<intersection>509 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>509,-100,509,-99</points>
<intersection>-100 1</intersection>
<intersection>-99 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>509,-99,534,-99</points>
<connection>
<GID>729</GID>
<name>IN_2</name></connection>
<connection>
<GID>746</GID>
<name>IN_2</name></connection>
<intersection>509 3</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591.5,-187.5,591.5,-182</points>
<intersection>-187.5 2</intersection>
<intersection>-182 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591.5,-182,624.5,-182</points>
<connection>
<GID>130</GID>
<name>IN_6</name></connection>
<intersection>591.5 0</intersection>
<intersection>604 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-187.5,591.5,-187.5</points>
<connection>
<GID>134</GID>
<name>OUT_3</name></connection>
<intersection>591.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>604,-182,604,-159</points>
<intersection>-182 1</intersection>
<intersection>-159 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>604,-159,624.5,-159</points>
<connection>
<GID>129</GID>
<name>IN_6</name></connection>
<intersection>604 3</intersection></hsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,-108.5,509.5,-101</points>
<intersection>-108.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,-108.5,534,-108.5</points>
<connection>
<GID>730</GID>
<name>IN_2</name></connection>
<connection>
<GID>747</GID>
<name>IN_2</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-101,509.5,-101</points>
<connection>
<GID>689</GID>
<name>OUT_4</name></connection>
<intersection>509.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592,-188.5,592,-184</points>
<intersection>-188.5 2</intersection>
<intersection>-184 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592,-184,624.5,-184</points>
<connection>
<GID>130</GID>
<name>IN_4</name></connection>
<intersection>592 0</intersection>
<intersection>605 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>588.5,-188.5,592,-188.5</points>
<connection>
<GID>134</GID>
<name>OUT_2</name></connection>
<intersection>592 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>605,-184,605,-161</points>
<intersection>-184 1</intersection>
<intersection>-161 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>605,-161,624.5,-161</points>
<connection>
<GID>129</GID>
<name>IN_4</name></connection>
<intersection>605 3</intersection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510,-119.5,510,-102</points>
<intersection>-119.5 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510,-119.5,534,-119.5</points>
<connection>
<GID>731</GID>
<name>IN_2</name></connection>
<connection>
<GID>748</GID>
<name>IN_2</name></connection>
<intersection>510 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-102,510,-102</points>
<connection>
<GID>689</GID>
<name>OUT_3</name></connection>
<intersection>510 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510.5,-130.5,510.5,-103</points>
<intersection>-130.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,-130.5,534,-130.5</points>
<connection>
<GID>732</GID>
<name>IN_2</name></connection>
<connection>
<GID>749</GID>
<name>IN_2</name></connection>
<intersection>510.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-103,510.5,-103</points>
<connection>
<GID>689</GID>
<name>OUT_2</name></connection>
<intersection>510.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511,-141,511,-104</points>
<intersection>-141 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,-104,511,-104</points>
<connection>
<GID>689</GID>
<name>OUT_1</name></connection>
<intersection>511 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>511,-141,534,-141</points>
<connection>
<GID>733</GID>
<name>IN_2</name></connection>
<connection>
<GID>750</GID>
<name>IN_2</name></connection>
<intersection>511 0</intersection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-152,511.5,-105</points>
<intersection>-152 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511.5,-152,534,-152</points>
<connection>
<GID>734</GID>
<name>IN_2</name></connection>
<connection>
<GID>751</GID>
<name>IN_2</name></connection>
<intersection>511.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-105,511.5,-105</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,-111.5,512.5,-79</points>
<intersection>-111.5 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512.5,-79,534,-79</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<connection>
<GID>744</GID>
<name>IN_1</name></connection>
<intersection>512.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-111.5,512.5,-111.5</points>
<connection>
<GID>725</GID>
<name>OUT_7</name></connection>
<intersection>512.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,-112.5,513,-90</points>
<intersection>-112.5 2</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513,-90,534,-90</points>
<connection>
<GID>728</GID>
<name>IN_1</name></connection>
<connection>
<GID>745</GID>
<name>IN_1</name></connection>
<intersection>513 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-112.5,513,-112.5</points>
<connection>
<GID>725</GID>
<name>OUT_6</name></connection>
<intersection>513 0</intersection></hsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513.5,-113.5,513.5,-101</points>
<intersection>-113.5 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>513.5,-101,534,-101</points>
<connection>
<GID>746</GID>
<name>IN_1</name></connection>
<connection>
<GID>729</GID>
<name>IN_1</name></connection>
<intersection>513.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-113.5,513.5,-113.5</points>
<connection>
<GID>725</GID>
<name>OUT_5</name></connection>
<intersection>513.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-114.5,514,-110.5</points>
<intersection>-114.5 2</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-110.5,534,-110.5</points>
<connection>
<GID>730</GID>
<name>IN_1</name></connection>
<connection>
<GID>747</GID>
<name>IN_1</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-114.5,514,-114.5</points>
<connection>
<GID>725</GID>
<name>OUT_4</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,-121.5,514.5,-115.5</points>
<intersection>-121.5 1</intersection>
<intersection>-115.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514.5,-121.5,534,-121.5</points>
<connection>
<GID>731</GID>
<name>IN_1</name></connection>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-115.5,514.5,-115.5</points>
<connection>
<GID>725</GID>
<name>OUT_3</name></connection>
<intersection>514.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515,-132.5,515,-116.5</points>
<intersection>-132.5 1</intersection>
<intersection>-116.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515,-132.5,534,-132.5</points>
<connection>
<GID>732</GID>
<name>IN_1</name></connection>
<connection>
<GID>749</GID>
<name>IN_1</name></connection>
<intersection>515 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,-116.5,515,-116.5</points>
<connection>
<GID>725</GID>
<name>OUT_2</name></connection>
<intersection>515 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>319.289,532.775,402.711,489.75</PageViewport>
<gate>
<ID>152</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>381,523.5</position>
<input>
<ID>IN_0</ID>930 </input>
<input>
<ID>IN_1</ID>922 </input>
<input>
<ID>IN_10</ID>925 </input>
<input>
<ID>IN_11</ID>917 </input>
<input>
<ID>IN_12</ID>924 </input>
<input>
<ID>IN_13</ID>916 </input>
<input>
<ID>IN_14</ID>923 </input>
<input>
<ID>IN_15</ID>915 </input>
<input>
<ID>IN_2</ID>929 </input>
<input>
<ID>IN_3</ID>921 </input>
<input>
<ID>IN_4</ID>928 </input>
<input>
<ID>IN_5</ID>920 </input>
<input>
<ID>IN_6</ID>927 </input>
<input>
<ID>IN_7</ID>919 </input>
<input>
<ID>IN_8</ID>926 </input>
<input>
<ID>IN_9</ID>918 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>154</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>381,500.5</position>
<input>
<ID>IN_0</ID>930 </input>
<input>
<ID>IN_1</ID>922 </input>
<input>
<ID>IN_10</ID>925 </input>
<input>
<ID>IN_11</ID>917 </input>
<input>
<ID>IN_12</ID>924 </input>
<input>
<ID>IN_13</ID>916 </input>
<input>
<ID>IN_14</ID>923 </input>
<input>
<ID>IN_15</ID>915 </input>
<input>
<ID>IN_2</ID>929 </input>
<input>
<ID>IN_3</ID>921 </input>
<input>
<ID>IN_4</ID>928 </input>
<input>
<ID>IN_5</ID>920 </input>
<input>
<ID>IN_6</ID>927 </input>
<input>
<ID>IN_7</ID>919 </input>
<input>
<ID>IN_8</ID>926 </input>
<input>
<ID>IN_9</ID>918 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>155</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>341,525.5</position>
<output>
<ID>OUT_0</ID>922 </output>
<output>
<ID>OUT_1</ID>921 </output>
<output>
<ID>OUT_2</ID>920 </output>
<output>
<ID>OUT_3</ID>919 </output>
<output>
<ID>OUT_4</ID>918 </output>
<output>
<ID>OUT_5</ID>917 </output>
<output>
<ID>OUT_6</ID>916 </output>
<output>
<ID>OUT_7</ID>915 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>156</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>341,494</position>
<input>
<ID>ENABLE_0</ID>931 </input>
<output>
<ID>OUT_0</ID>930 </output>
<output>
<ID>OUT_1</ID>929 </output>
<output>
<ID>OUT_2</ID>928 </output>
<output>
<ID>OUT_3</ID>927 </output>
<output>
<ID>OUT_4</ID>926 </output>
<output>
<ID>OUT_5</ID>925 </output>
<output>
<ID>OUT_6</ID>924 </output>
<output>
<ID>OUT_7</ID>923 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>158</ID>
<type>EE_VDD</type>
<position>341,509</position>
<output>
<ID>OUT_0</ID>931 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,529,351.5,531</points>
<intersection>529 2</intersection>
<intersection>531 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,531,379,531</points>
<connection>
<GID>152</GID>
<name>IN_15</name></connection>
<intersection>351.5 0</intersection>
<intersection>354 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,529,351.5,529</points>
<connection>
<GID>155</GID>
<name>OUT_7</name></connection>
<intersection>351.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>354,508,354,531</points>
<intersection>508 4</intersection>
<intersection>531 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354,508,379,508</points>
<connection>
<GID>154</GID>
<name>IN_15</name></connection>
<intersection>354 3</intersection></hsegment></shape></wire>
<wire>
<ID>916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,528,352,529</points>
<intersection>528 2</intersection>
<intersection>529 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,529,379,529</points>
<connection>
<GID>152</GID>
<name>IN_13</name></connection>
<intersection>352 0</intersection>
<intersection>355 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,528,352,528</points>
<connection>
<GID>155</GID>
<name>OUT_6</name></connection>
<intersection>352 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>355,506,355,529</points>
<intersection>506 4</intersection>
<intersection>529 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355,506,379,506</points>
<connection>
<GID>154</GID>
<name>IN_13</name></connection>
<intersection>355 3</intersection></hsegment></shape></wire>
<wire>
<ID>917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343,527,379,527</points>
<connection>
<GID>155</GID>
<name>OUT_5</name></connection>
<connection>
<GID>152</GID>
<name>IN_11</name></connection>
<intersection>357 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>357,504,357,527</points>
<intersection>504 3</intersection>
<intersection>527 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>357,504,379,504</points>
<connection>
<GID>154</GID>
<name>IN_11</name></connection>
<intersection>357 2</intersection></hsegment></shape></wire>
<wire>
<ID>918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351.5,525,351.5,526</points>
<intersection>525 1</intersection>
<intersection>526 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351.5,525,379,525</points>
<connection>
<GID>152</GID>
<name>IN_9</name></connection>
<intersection>351.5 0</intersection>
<intersection>357 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,526,351.5,526</points>
<connection>
<GID>155</GID>
<name>OUT_4</name></connection>
<intersection>351.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>357,502,357,525</points>
<intersection>502 4</intersection>
<intersection>525 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>357,502,379,502</points>
<connection>
<GID>154</GID>
<name>IN_9</name></connection>
<intersection>357 3</intersection></hsegment></shape></wire>
<wire>
<ID>919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,523,351,525</points>
<intersection>523 1</intersection>
<intersection>525 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,523,379,523</points>
<connection>
<GID>152</GID>
<name>IN_7</name></connection>
<intersection>351 0</intersection>
<intersection>358 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,525,351,525</points>
<connection>
<GID>155</GID>
<name>OUT_3</name></connection>
<intersection>351 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>358,500,358,523</points>
<intersection>500 4</intersection>
<intersection>523 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>358,500,379,500</points>
<connection>
<GID>154</GID>
<name>IN_7</name></connection>
<intersection>358 3</intersection></hsegment></shape></wire>
<wire>
<ID>920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350.5,521,350.5,524</points>
<intersection>521 1</intersection>
<intersection>524 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350.5,521,379,521</points>
<connection>
<GID>152</GID>
<name>IN_5</name></connection>
<intersection>350.5 0</intersection>
<intersection>359 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,524,350.5,524</points>
<connection>
<GID>155</GID>
<name>OUT_2</name></connection>
<intersection>350.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>359,498,359,521</points>
<intersection>498 4</intersection>
<intersection>521 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>359,498,379,498</points>
<connection>
<GID>154</GID>
<name>IN_5</name></connection>
<intersection>359 3</intersection></hsegment></shape></wire>
<wire>
<ID>921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,519,350,523</points>
<intersection>519 1</intersection>
<intersection>523 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,519,379,519</points>
<connection>
<GID>152</GID>
<name>IN_3</name></connection>
<intersection>350 0</intersection>
<intersection>360 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,523,350,523</points>
<connection>
<GID>155</GID>
<name>OUT_1</name></connection>
<intersection>350 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>360,496,360,519</points>
<intersection>496 4</intersection>
<intersection>519 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>360,496,379,496</points>
<connection>
<GID>154</GID>
<name>IN_3</name></connection>
<intersection>360 3</intersection></hsegment></shape></wire>
<wire>
<ID>922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,517,349.5,522</points>
<intersection>517 1</intersection>
<intersection>522 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349.5,517,379,517</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>349.5 0</intersection>
<intersection>361 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,522,349.5,522</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>361,494,361,517</points>
<intersection>494 4</intersection>
<intersection>517 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>361,494,379,494</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>361 3</intersection></hsegment></shape></wire>
<wire>
<ID>923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,497.5,344,507</points>
<intersection>497.5 2</intersection>
<intersection>507 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,507,379,507</points>
<connection>
<GID>154</GID>
<name>IN_14</name></connection>
<intersection>344 0</intersection>
<intersection>354.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,497.5,344,497.5</points>
<connection>
<GID>156</GID>
<name>OUT_7</name></connection>
<intersection>344 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>354.5,507,354.5,530</points>
<intersection>507 1</intersection>
<intersection>530 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>354.5,530,379,530</points>
<connection>
<GID>152</GID>
<name>IN_14</name></connection>
<intersection>354.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>924</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,496.5,344.5,505</points>
<intersection>496.5 2</intersection>
<intersection>505 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,505,379,505</points>
<connection>
<GID>154</GID>
<name>IN_12</name></connection>
<intersection>344.5 0</intersection>
<intersection>355.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,496.5,344.5,496.5</points>
<connection>
<GID>156</GID>
<name>OUT_6</name></connection>
<intersection>344.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>355.5,505,355.5,528</points>
<intersection>505 1</intersection>
<intersection>528 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>355.5,528,379,528</points>
<connection>
<GID>152</GID>
<name>IN_12</name></connection>
<intersection>355.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>925</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345,495.5,345,503</points>
<intersection>495.5 2</intersection>
<intersection>503 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345,503,379,503</points>
<connection>
<GID>154</GID>
<name>IN_10</name></connection>
<intersection>345 0</intersection>
<intersection>356.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,495.5,345,495.5</points>
<connection>
<GID>156</GID>
<name>OUT_5</name></connection>
<intersection>345 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>356.5,503,356.5,526</points>
<intersection>503 1</intersection>
<intersection>526 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>356.5,526,379,526</points>
<connection>
<GID>152</GID>
<name>IN_10</name></connection>
<intersection>356.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>926</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345.5,494.5,345.5,501</points>
<intersection>494.5 2</intersection>
<intersection>501 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345.5,501,379,501</points>
<connection>
<GID>154</GID>
<name>IN_8</name></connection>
<intersection>345.5 0</intersection>
<intersection>357.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,494.5,345.5,494.5</points>
<connection>
<GID>156</GID>
<name>OUT_4</name></connection>
<intersection>345.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>357.5,501,357.5,524</points>
<intersection>501 1</intersection>
<intersection>524 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>357.5,524,379,524</points>
<connection>
<GID>152</GID>
<name>IN_8</name></connection>
<intersection>357.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>927</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346,493.5,346,499</points>
<intersection>493.5 2</intersection>
<intersection>499 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346,499,379,499</points>
<connection>
<GID>154</GID>
<name>IN_6</name></connection>
<intersection>346 0</intersection>
<intersection>358.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,493.5,346,493.5</points>
<connection>
<GID>156</GID>
<name>OUT_3</name></connection>
<intersection>346 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>358.5,499,358.5,522</points>
<intersection>499 1</intersection>
<intersection>522 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>358.5,522,379,522</points>
<connection>
<GID>152</GID>
<name>IN_6</name></connection>
<intersection>358.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>928</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346.5,492.5,346.5,497</points>
<intersection>492.5 2</intersection>
<intersection>497 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346.5,497,379,497</points>
<connection>
<GID>154</GID>
<name>IN_4</name></connection>
<intersection>346.5 0</intersection>
<intersection>359.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,492.5,346.5,492.5</points>
<connection>
<GID>156</GID>
<name>OUT_2</name></connection>
<intersection>346.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>359.5,497,359.5,520</points>
<intersection>497 1</intersection>
<intersection>520 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>359.5,520,379,520</points>
<connection>
<GID>152</GID>
<name>IN_4</name></connection>
<intersection>359.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>929</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,491.5,347,495</points>
<intersection>491.5 2</intersection>
<intersection>495 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,495,379,495</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<intersection>347 0</intersection>
<intersection>360.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,491.5,347,491.5</points>
<connection>
<GID>156</GID>
<name>OUT_1</name></connection>
<intersection>347 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>360.5,495,360.5,518</points>
<intersection>495 1</intersection>
<intersection>518 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>360.5,518,379,518</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>360.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347.5,490.5,347.5,493</points>
<intersection>490.5 2</intersection>
<intersection>493 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347.5,493,379,493</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>347.5 0</intersection>
<intersection>361.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343,490.5,347.5,490.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<intersection>347.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>361.5,493,361.5,516</points>
<intersection>493 1</intersection>
<intersection>516 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>361.5,516,379,516</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>361.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>341,499,341,508</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>-10.866,748.48,1767.13,-168.52</PageViewport></page 8>
<page 9>
<PageViewport>-10.866,748.48,1767.13,-168.52</PageViewport></page 9></circuit>