<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-87.8065,-184.572,281.419,-344.46</PageViewport>
<gate>
<ID>3</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>101,-297</position>
<input>
<ID>ENABLE_0</ID>83 </input>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_4</ID>55 </input>
<input>
<ID>IN_5</ID>56 </input>
<input>
<ID>IN_6</ID>57 </input>
<input>
<ID>IN_7</ID>58 </input>
<output>
<ID>OUT_0</ID>82 </output>
<output>
<ID>OUT_1</ID>81 </output>
<output>
<ID>OUT_2</ID>80 </output>
<output>
<ID>OUT_3</ID>79 </output>
<output>
<ID>OUT_4</ID>78 </output>
<output>
<ID>OUT_5</ID>77 </output>
<output>
<ID>OUT_6</ID>76 </output>
<output>
<ID>OUT_7</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_MUX_4x1</type>
<position>54,-294.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>63 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_MUX_4x1</type>
<position>54,-305</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>64 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_MUX_4x1</type>
<position>54,-316.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>65 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_MUX_4x1</type>
<position>54,-327.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>66 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_MUX_4x1</type>
<position>53.5,-272</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>61 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_MUX_4x1</type>
<position>54,-262</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>60 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_MUX_4x1</type>
<position>53.5,-251</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>59 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>96.5,-286</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Gate.PC</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>53,-237</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MUX0.PC</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>52,-240.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MUX1.PC</lparam></gate>
<gate>
<ID>14</ID>
<type>BM_ROM_16x16</type>
<position>193,-265</position>
<input>
<ID>ADDRESS_0</ID>96 </input>
<input>
<ID>ADDRESS_1</ID>97 </input>
<input>
<ID>ADDRESS_2</ID>98 </input>
<input>
<ID>ADDRESS_3</ID>99 </input>
<output>
<ID>DATA_OUT_10</ID>109 </output>
<output>
<ID>DATA_OUT_11</ID>94 </output>
<output>
<ID>DATA_OUT_12</ID>93 </output>
<output>
<ID>DATA_OUT_13</ID>92 </output>
<output>
<ID>DATA_OUT_14</ID>91 </output>
<output>
<ID>DATA_OUT_15</ID>90 </output>
<output>
<ID>DATA_OUT_8</ID>95 </output>
<output>
<ID>DATA_OUT_9</ID>108 </output>
<input>
<ID>ENABLE_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 16</lparam>
<lparam>DATA_BITS 16</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>201,-286</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R.MEM</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>201,-290</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W.MEM</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>201,-294.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD.PC</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>201,-299</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Gate.PC</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>201,-303</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MUX0.PC</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>201,-306.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MUX1.PC</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>200.5,-310.5</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD.IR</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>82.5,-326.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>6.5,-370</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_TO</type>
<position>201,-283</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>205,-258</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>DD_KEYPAD_HEX</type>
<position>170,-269.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<output>
<ID>OUT_1</ID>97 </output>
<output>
<ID>OUT_2</ID>98 </output>
<output>
<ID>OUT_3</ID>99 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>DD_KEYPAD_HEX</type>
<position>3,-232</position>
<output>
<ID>OUT_0</ID>104 </output>
<output>
<ID>OUT_1</ID>105 </output>
<output>
<ID>OUT_2</ID>106 </output>
<output>
<ID>OUT_3</ID>107 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>28</ID>
<type>DD_KEYPAD_HEX</type>
<position>2.5,-245.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<output>
<ID>OUT_1</ID>101 </output>
<output>
<ID>OUT_2</ID>102 </output>
<output>
<ID>OUT_3</ID>103 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 14</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_RAM_8x8</type>
<position>86,-386.5</position>
<input>
<ID>ADDRESS_0</ID>36 </input>
<input>
<ID>ADDRESS_1</ID>35 </input>
<input>
<ID>ADDRESS_2</ID>34 </input>
<input>
<ID>ADDRESS_3</ID>33 </input>
<input>
<ID>ADDRESS_4</ID>32 </input>
<input>
<ID>ADDRESS_5</ID>31 </input>
<input>
<ID>ADDRESS_6</ID>30 </input>
<input>
<ID>ADDRESS_7</ID>29 </input>
<input>
<ID>DATA_IN_0</ID>8 </input>
<input>
<ID>DATA_IN_1</ID>7 </input>
<input>
<ID>DATA_IN_2</ID>6 </input>
<input>
<ID>DATA_IN_3</ID>5 </input>
<input>
<ID>DATA_IN_4</ID>4 </input>
<input>
<ID>DATA_IN_5</ID>3 </input>
<input>
<ID>DATA_IN_6</ID>2 </input>
<input>
<ID>DATA_IN_7</ID>1 </input>
<output>
<ID>DATA_OUT_0</ID>8 </output>
<output>
<ID>DATA_OUT_1</ID>7 </output>
<output>
<ID>DATA_OUT_2</ID>6 </output>
<output>
<ID>DATA_OUT_3</ID>5 </output>
<output>
<ID>DATA_OUT_4</ID>4 </output>
<output>
<ID>DATA_OUT_5</ID>3 </output>
<output>
<ID>DATA_OUT_6</ID>2 </output>
<output>
<ID>DATA_OUT_7</ID>1 </output>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>write_clock</ID>11 </input>
<input>
<ID>write_enable</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>30</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>93.5,-400.5</position>
<input>
<ID>ENABLE_0</ID>28 </input>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>3 </input>
<input>
<ID>IN_6</ID>2 </input>
<input>
<ID>IN_7</ID>1 </input>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>25 </output>
<output>
<ID>OUT_2</ID>24 </output>
<output>
<ID>OUT_3</ID>23 </output>
<output>
<ID>OUT_4</ID>22 </output>
<output>
<ID>OUT_5</ID>21 </output>
<output>
<ID>OUT_6</ID>20 </output>
<output>
<ID>OUT_7</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>31</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>80,-400.5</position>
<input>
<ID>ENABLE_0</ID>27 </input>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>15 </input>
<input>
<ID>IN_4</ID>12 </input>
<input>
<ID>IN_5</ID>14 </input>
<input>
<ID>IN_6</ID>13 </input>
<input>
<ID>IN_7</ID>9 </input>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>7 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>5 </output>
<output>
<ID>OUT_4</ID>4 </output>
<output>
<ID>OUT_5</ID>3 </output>
<output>
<ID>OUT_6</ID>2 </output>
<output>
<ID>OUT_7</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>32</ID>
<type>BB_CLOCK</type>
<position>170,-248.5</position>
<output>
<ID>CLK</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 4</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>62.5,-393</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>62.5,-395</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>180.5,-249</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>103.5,-385</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>62.5,-397</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>62.5,-399</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>62.5,-401.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>62.5,-404</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>62.5,-406</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>62.5,-408.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>101,-394</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>101,-396.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>101,-398.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>101,-400.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>101,-403</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>101,-405</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>101,-407.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>101,-410</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>63,-381</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID W.MEM</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>63,-378.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R.MEM</lparam></gate>
<gate>
<ID>53</ID>
<type>DA_FROM</type>
<position>48.5,-382</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>48.5,-384</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>48.5,-386</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>48.5,-388</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>48.5,-390.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>48.5,-393</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>48.5,-395</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>48.5,-397.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_REGISTER8</type>
<position>84.5,-311</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>61 </input>
<input>
<ID>IN_6</ID>60 </input>
<input>
<ID>IN_7</ID>59 </input>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>52 </output>
<output>
<ID>OUT_2</ID>53 </output>
<output>
<ID>OUT_3</ID>54 </output>
<output>
<ID>OUT_4</ID>55 </output>
<output>
<ID>OUT_5</ID>56 </output>
<output>
<ID>OUT_6</ID>57 </output>
<output>
<ID>OUT_7</ID>58 </output>
<input>
<ID>clear</ID>87 </input>
<input>
<ID>clock</ID>45 </input>
<input>
<ID>load</ID>86 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 254</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_REGISTER8</type>
<position>9.5,-356.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<input>
<ID>IN_4</ID>40 </input>
<input>
<ID>IN_5</ID>39 </input>
<input>
<ID>IN_6</ID>38 </input>
<input>
<ID>IN_7</ID>37 </input>
<input>
<ID>clear</ID>88 </input>
<input>
<ID>clock</ID>46 </input>
<input>
<ID>load</ID>47 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 204</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>6.5,-362</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>84,-317.5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-6,-349</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>-6,-351</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>-6,-353</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>-6,-355</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>-6,-357.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>-6,-360</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>-6,-362</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>-6,-364.5</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>110.5,-288</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>110.5,-290.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>110.5,-292.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>110.5,-294.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>110.5,-297</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>110.5,-299</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>110.5,-301.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>110.5,-304</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>78.5,-322</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>5,-367</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>79,-298</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD.PC</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-9.5,-345</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD.IR</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_FULLADDER_4BIT</type>
<position>138,-329.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_B_0</ID>50 </input>
<input>
<ID>IN_B_1</ID>49 </input>
<input>
<ID>IN_B_2</ID>49 </input>
<input>
<ID>IN_B_3</ID>49 </input>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>68 </output>
<output>
<ID>OUT_2</ID>69 </output>
<output>
<ID>OUT_3</ID>70 </output>
<output>
<ID>carry_out</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_FULLADDER_4BIT</type>
<position>119.5,-329.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>58 </input>
<input>
<ID>IN_B_0</ID>49 </input>
<input>
<ID>IN_B_1</ID>49 </input>
<input>
<ID>IN_B_2</ID>49 </input>
<input>
<ID>IN_B_3</ID>49 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<input>
<ID>carry_in</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>87</ID>
<type>FF_GND</type>
<position>120.5,-317.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>EE_VDD</type>
<position>143,-314.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_MUX_4x1</type>
<position>54,-284</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>62 </output>
<input>
<ID>SEL_0</ID>84 </input>
<input>
<ID>SEL_1</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-397,82.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_7</name></connection>
<intersection>-397 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-397,91.5,-397</points>
<connection>
<GID>30</GID>
<name>IN_7</name></connection>
<connection>
<GID>31</GID>
<name>OUT_7</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-398,83.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_6</name></connection>
<intersection>-398 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-398,91.5,-398</points>
<connection>
<GID>30</GID>
<name>IN_6</name></connection>
<connection>
<GID>31</GID>
<name>OUT_6</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-399,84.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_5</name></connection>
<intersection>-399 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-399,91.5,-399</points>
<connection>
<GID>30</GID>
<name>IN_5</name></connection>
<connection>
<GID>31</GID>
<name>OUT_5</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-400,85.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_4</name></connection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-400,91.5,-400</points>
<connection>
<GID>30</GID>
<name>IN_4</name></connection>
<connection>
<GID>31</GID>
<name>OUT_4</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-401,86.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_3</name></connection>
<intersection>-401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-401,91.5,-401</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-402,87.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_2</name></connection>
<intersection>-402 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-402,91.5,-402</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-403,88.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_1</name></connection>
<intersection>-403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-403,91.5,-403</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-404,89.5,-393.5</points>
<connection>
<GID>29</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>DATA_IN_0</name></connection>
<intersection>-404 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-404,91.5,-404</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-393,78,-393</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>78 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78,-397,78,-393</points>
<connection>
<GID>31</GID>
<name>IN_7</name></connection>
<intersection>-393 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>174,-248.5,178.5,-248.5</points>
<connection>
<GID>32</GID>
<name>CLK</name></connection>
<intersection>178.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>178.5,-249,178.5,-248.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>-248.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91,-385,105.5,-385</points>
<connection>
<GID>29</GID>
<name>write_clock</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-400,77.5,-399</points>
<intersection>-400 1</intersection>
<intersection>-399 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-400,78,-400</points>
<connection>
<GID>31</GID>
<name>IN_4</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-399,77.5,-399</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-398,77,-395</points>
<intersection>-398 1</intersection>
<intersection>-395 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-398,78,-398</points>
<connection>
<GID>31</GID>
<name>IN_6</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-395,77,-395</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-399,77.5,-397</points>
<intersection>-399 1</intersection>
<intersection>-397 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-399,78,-399</points>
<connection>
<GID>31</GID>
<name>IN_5</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-397,77.5,-397</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-401.5,77.5,-401</points>
<intersection>-401.5 2</intersection>
<intersection>-401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-401,78,-401</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-401.5,77.5,-401.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-408.5,77.5,-404</points>
<intersection>-408.5 2</intersection>
<intersection>-404 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-404,78,-404</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-408.5,77.5,-408.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-404,77.5,-402</points>
<intersection>-404 2</intersection>
<intersection>-402 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-402,78,-402</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-404,77.5,-404</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-406,77.5,-403</points>
<intersection>-406 2</intersection>
<intersection>-403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-403,78,-403</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-406,77.5,-406</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-397,97,-394</points>
<intersection>-397 2</intersection>
<intersection>-394 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-394,99,-394</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-397,97,-397</points>
<connection>
<GID>30</GID>
<name>OUT_7</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-398,97,-396.5</points>
<intersection>-398 1</intersection>
<intersection>-396.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-398,97,-398</points>
<connection>
<GID>30</GID>
<name>OUT_6</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-396.5,99,-396.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-399,97,-398.5</points>
<intersection>-399 1</intersection>
<intersection>-398.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-399,97,-399</points>
<connection>
<GID>30</GID>
<name>OUT_5</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-398.5,99,-398.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-400.5,97,-400</points>
<intersection>-400.5 2</intersection>
<intersection>-400 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-400,97,-400</points>
<connection>
<GID>30</GID>
<name>OUT_4</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-400.5,99,-400.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-403,97,-401</points>
<intersection>-403 2</intersection>
<intersection>-401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-401,97,-401</points>
<connection>
<GID>30</GID>
<name>OUT_3</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-403,99,-403</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-405,97,-402</points>
<intersection>-405 2</intersection>
<intersection>-402 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-402,97,-402</points>
<connection>
<GID>30</GID>
<name>OUT_2</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-405,99,-405</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-407.5,97,-403</points>
<intersection>-407.5 2</intersection>
<intersection>-403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-403,97,-403</points>
<connection>
<GID>30</GID>
<name>OUT_1</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-407.5,99,-407.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-410,97,-404</points>
<intersection>-410 2</intersection>
<intersection>-404 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-404,97,-404</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-410,99,-410</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-379,91.5,-379</points>
<intersection>65 7</intersection>
<intersection>91 10</intersection>
<intersection>91.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-395.5,91.5,-379</points>
<intersection>-395.5 4</intersection>
<intersection>-379 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>80,-395.5,91.5,-395.5</points>
<connection>
<GID>31</GID>
<name>ENABLE_0</name></connection>
<intersection>91.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>65,-381,65,-379</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-379 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>91,-386,91,-379</points>
<connection>
<GID>29</GID>
<name>write_enable</name></connection>
<intersection>-379 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65,-378.5,93.5,-378.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>91 3</intersection>
<intersection>93.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91,-387,91,-378.5</points>
<connection>
<GID>29</GID>
<name>ENABLE_0</name></connection>
<intersection>-378.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>93.5,-395.5,93.5,-378.5</points>
<connection>
<GID>30</GID>
<name>ENABLE_0</name></connection>
<intersection>-378.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-383,65.5,-382</points>
<intersection>-383 1</intersection>
<intersection>-382 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-383,81,-383</points>
<connection>
<GID>29</GID>
<name>ADDRESS_7</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-382,65.5,-382</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-384,81,-384</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-386,65.5,-385</points>
<intersection>-386 2</intersection>
<intersection>-385 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-385,81,-385</points>
<connection>
<GID>29</GID>
<name>ADDRESS_5</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-386,65.5,-386</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-388,65.5,-386</points>
<intersection>-388 2</intersection>
<intersection>-386 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-386,81,-386</points>
<connection>
<GID>29</GID>
<name>ADDRESS_4</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-388,65.5,-388</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-390.5,65.5,-387</points>
<intersection>-390.5 2</intersection>
<intersection>-387 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-387,81,-387</points>
<connection>
<GID>29</GID>
<name>ADDRESS_3</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-390.5,65.5,-390.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-393,65.5,-388</points>
<intersection>-393 2</intersection>
<intersection>-388 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-388,81,-388</points>
<connection>
<GID>29</GID>
<name>ADDRESS_2</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-393,65.5,-393</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-395,65.5,-389</points>
<intersection>-395 2</intersection>
<intersection>-389 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-389,81,-389</points>
<connection>
<GID>29</GID>
<name>ADDRESS_1</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-395,65.5,-395</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-397.5,65.5,-390</points>
<intersection>-397.5 2</intersection>
<intersection>-390 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-390,81,-390</points>
<connection>
<GID>29</GID>
<name>ADDRESS_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-397.5,65.5,-397.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-352.5,0.5,-349</points>
<intersection>-352.5 1</intersection>
<intersection>-349 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-352.5,5.5,-352.5</points>
<connection>
<GID>62</GID>
<name>IN_7</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-349,0.5,-349</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-353.5,0.5,-351</points>
<intersection>-353.5 1</intersection>
<intersection>-351 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-353.5,5.5,-353.5</points>
<connection>
<GID>62</GID>
<name>IN_6</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-351,0.5,-351</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-354.5,0.5,-353</points>
<intersection>-354.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-354.5,5.5,-354.5</points>
<connection>
<GID>62</GID>
<name>IN_5</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-353,0.5,-353</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-355.5,0.5,-355</points>
<intersection>-355.5 1</intersection>
<intersection>-355 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-355.5,5.5,-355.5</points>
<connection>
<GID>62</GID>
<name>IN_4</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-355,0.5,-355</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-357.5,0.5,-356.5</points>
<intersection>-357.5 2</intersection>
<intersection>-356.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-356.5,5.5,-356.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-357.5,0.5,-357.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-360,0.5,-357.5</points>
<intersection>-360 2</intersection>
<intersection>-357.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-357.5,5.5,-357.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-360,0.5,-360</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-362,0.5,-358.5</points>
<intersection>-362 2</intersection>
<intersection>-358.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-358.5,5.5,-358.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-362,0.5,-362</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-364.5,0.5,-359.5</points>
<intersection>-364.5 2</intersection>
<intersection>-359.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-359.5,5.5,-359.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-364.5,0.5,-364.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-322,83.5,-316</points>
<connection>
<GID>61</GID>
<name>clock</name></connection>
<intersection>-322 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-322,83.5,-322</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-367,8.5,-361.5</points>
<connection>
<GID>62</GID>
<name>clock</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-367,8.5,-367</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-350.5,8.5,-345</points>
<connection>
<GID>62</GID>
<name>load</name></connection>
<intersection>-345 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-345,8.5,-345</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-328.5,130,-328.5</points>
<connection>
<GID>86</GID>
<name>carry_in</name></connection>
<connection>
<GID>85</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-325.5,121.5,-317.5</points>
<connection>
<GID>86</GID>
<name>IN_B_3</name></connection>
<intersection>-319 4</intersection>
<intersection>-317.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>122.5,-317.5,122.5,-316.5</points>
<intersection>-317.5 2</intersection>
<intersection>-316.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-317.5,122.5,-317.5</points>
<intersection>121.5 0</intersection>
<intersection>122.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>120.5,-316.5,122.5,-316.5</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>122.5 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>121.5,-319,142,-319</points>
<intersection>121.5 0</intersection>
<intersection>122.5 16</intersection>
<intersection>123.5 15</intersection>
<intersection>124.5 14</intersection>
<intersection>140 13</intersection>
<intersection>141 12</intersection>
<intersection>142 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>142,-325.5,142,-319</points>
<connection>
<GID>85</GID>
<name>IN_B_1</name></connection>
<intersection>-319 4</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>141,-325.5,141,-319</points>
<connection>
<GID>85</GID>
<name>IN_B_2</name></connection>
<intersection>-319 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>140,-325.5,140,-319</points>
<connection>
<GID>85</GID>
<name>IN_B_3</name></connection>
<intersection>-319 4</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>124.5,-325.5,124.5,-319</points>
<connection>
<GID>86</GID>
<name>IN_B_0</name></connection>
<intersection>-319 4</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>123.5,-325.5,123.5,-319</points>
<connection>
<GID>86</GID>
<name>IN_B_1</name></connection>
<intersection>-319 4</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>122.5,-325.5,122.5,-319</points>
<connection>
<GID>86</GID>
<name>IN_B_2</name></connection>
<intersection>-319 4</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-325.5,143,-315.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-325.5,136,-314</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-314 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-314,136,-314</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>98 2</intersection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-314,98,-300.5</points>
<intersection>-314 1</intersection>
<intersection>-300.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>98,-300.5,99,-300.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>98 2</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-325.5,135,-313</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-313,135,-313</points>
<connection>
<GID>61</GID>
<name>OUT_1</name></connection>
<intersection>97 2</intersection>
<intersection>135 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>97,-313,97,-299.5</points>
<intersection>-313 1</intersection>
<intersection>-299.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>97,-299.5,99,-299.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>97 2</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-325.5,134,-312</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>-312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-312,134,-312</points>
<connection>
<GID>61</GID>
<name>OUT_2</name></connection>
<intersection>96 2</intersection>
<intersection>134 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96,-312,96,-298.5</points>
<intersection>-312 1</intersection>
<intersection>-298.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>96,-298.5,99,-298.5</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>96 2</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-325.5,133,-311</points>
<connection>
<GID>85</GID>
<name>IN_3</name></connection>
<intersection>-311 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-311,133,-311</points>
<connection>
<GID>61</GID>
<name>OUT_3</name></connection>
<intersection>95 2</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>95,-311,95,-297.5</points>
<intersection>-311 1</intersection>
<intersection>-297.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95,-297.5,99,-297.5</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>95 2</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-325.5,117.5,-310</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>-310 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-310,117.5,-310</points>
<connection>
<GID>61</GID>
<name>OUT_4</name></connection>
<intersection>94 2</intersection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>94,-310,94,-296.5</points>
<intersection>-310 1</intersection>
<intersection>-296.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>94,-296.5,99,-296.5</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>94 2</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-325.5,116.5,-309</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>-309 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-309,116.5,-309</points>
<connection>
<GID>61</GID>
<name>OUT_5</name></connection>
<intersection>92.5 2</intersection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>92.5,-309,92.5,-295.5</points>
<intersection>-309 1</intersection>
<intersection>-295.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>92.5,-295.5,99,-295.5</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>92.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-325.5,115.5,-308</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>-308 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-308,115.5,-308</points>
<connection>
<GID>61</GID>
<name>OUT_6</name></connection>
<intersection>91.5 2</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>91.5,-308,91.5,-294.5</points>
<intersection>-308 1</intersection>
<intersection>-294.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>91.5,-294.5,99,-294.5</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>91.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-325.5,114.5,-307</points>
<connection>
<GID>86</GID>
<name>IN_3</name></connection>
<intersection>-307 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-307,114.5,-307</points>
<connection>
<GID>61</GID>
<name>OUT_7</name></connection>
<intersection>90.5 2</intersection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>90.5,-307,90.5,-293.5</points>
<intersection>-307 1</intersection>
<intersection>-293.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>90.5,-293.5,99,-293.5</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>90.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-307,68.5,-251</points>
<intersection>-307 1</intersection>
<intersection>-251 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-307,80.5,-307</points>
<connection>
<GID>61</GID>
<name>IN_7</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-251,68.5,-251</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-308,68.5,-262</points>
<intersection>-308 1</intersection>
<intersection>-262 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-308,80.5,-308</points>
<connection>
<GID>61</GID>
<name>IN_6</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-262,68.5,-262</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-309,68.5,-272</points>
<intersection>-309 1</intersection>
<intersection>-272 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-309,80.5,-309</points>
<connection>
<GID>61</GID>
<name>IN_5</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-272,68.5,-272</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-310,68.5,-284</points>
<intersection>-310 1</intersection>
<intersection>-284 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-310,80.5,-310</points>
<connection>
<GID>61</GID>
<name>IN_4</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-284,68.5,-284</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-311,68.5,-294.5</points>
<intersection>-311 1</intersection>
<intersection>-294.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-311,80.5,-311</points>
<connection>
<GID>61</GID>
<name>IN_3</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-294.5,68.5,-294.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-312,68.5,-305</points>
<intersection>-312 1</intersection>
<intersection>-305 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-312,80.5,-312</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-305,68.5,-305</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-316.5,68.5,-313</points>
<intersection>-316.5 2</intersection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-313,80.5,-313</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-316.5,68.5,-316.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-327.5,68.5,-314</points>
<intersection>-327.5 2</intersection>
<intersection>-314 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-314,80.5,-314</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-327.5,68.5,-327.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-337,139.5,-333.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>-337 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-337,139.5,-337</points>
<intersection>51 2</intersection>
<intersection>139.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>51,-337,51,-330.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-337 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-339,138.5,-333.5</points>
<connection>
<GID>85</GID>
<name>OUT_1</name></connection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-339,138.5,-339</points>
<intersection>49.5 2</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>49.5,-339,49.5,-319.5</points>
<intersection>-339 1</intersection>
<intersection>-319.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49.5,-319.5,51,-319.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>49.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-342,137.5,-333.5</points>
<connection>
<GID>85</GID>
<name>OUT_2</name></connection>
<intersection>-342 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-342,137.5,-342</points>
<intersection>49 2</intersection>
<intersection>137.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>49,-342,49,-308</points>
<intersection>-342 1</intersection>
<intersection>-308 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49,-308,51,-308</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>49 2</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-340.5,136.5,-333.5</points>
<connection>
<GID>85</GID>
<name>OUT_3</name></connection>
<intersection>-340.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-340.5,136.5,-340.5</points>
<intersection>48 2</intersection>
<intersection>136.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48,-340.5,48,-297.5</points>
<intersection>-340.5 1</intersection>
<intersection>-297.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>48,-297.5,51,-297.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>48 2</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-343,121,-333.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-343 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-343,121,-343</points>
<intersection>45.5 2</intersection>
<intersection>121 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>45.5,-343,45.5,-287</points>
<intersection>-343 1</intersection>
<intersection>-287 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>45.5,-287,51,-287</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>45.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-345.5,120,-333.5</points>
<connection>
<GID>86</GID>
<name>OUT_1</name></connection>
<intersection>-345.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-345.5,120,-345.5</points>
<intersection>43.5 2</intersection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>43.5,-345.5,43.5,-275</points>
<intersection>-345.5 1</intersection>
<intersection>-275 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>43.5,-275,50.5,-275</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>43.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-348.5,119,-333.5</points>
<connection>
<GID>86</GID>
<name>OUT_2</name></connection>
<intersection>-348.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-348.5,119,-348.5</points>
<intersection>41.5 2</intersection>
<intersection>119 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>41.5,-348.5,41.5,-265</points>
<intersection>-348.5 1</intersection>
<intersection>-265 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-265,51,-265</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>41.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-351,118,-333.5</points>
<connection>
<GID>86</GID>
<name>OUT_3</name></connection>
<intersection>-351 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-351,118,-351</points>
<intersection>40.5 2</intersection>
<intersection>118 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>40.5,-351,40.5,-254</points>
<intersection>-351 1</intersection>
<intersection>-254 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40.5,-254,50.5,-254</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>40.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-293.5,105,-288</points>
<intersection>-293.5 2</intersection>
<intersection>-288 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-288,108.5,-288</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-293.5,105,-293.5</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-294.5,105,-290.5</points>
<intersection>-294.5 2</intersection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-290.5,108.5,-290.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-294.5,105,-294.5</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-295.5,105,-292.5</points>
<intersection>-295.5 2</intersection>
<intersection>-292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-292.5,108.5,-292.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-295.5,105,-295.5</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-296.5,105.5,-294.5</points>
<intersection>-296.5 1</intersection>
<intersection>-294.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-296.5,105.5,-296.5</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-294.5,108.5,-294.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-297.5,105.5,-297</points>
<intersection>-297.5 2</intersection>
<intersection>-297 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-297,108.5,-297</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-297.5,105.5,-297.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-299,105.5,-298.5</points>
<intersection>-299 1</intersection>
<intersection>-298.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-299,108.5,-299</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-298.5,105.5,-298.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-301.5,105.5,-299.5</points>
<intersection>-301.5 1</intersection>
<intersection>-299.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-301.5,108.5,-301.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-299.5,105.5,-299.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-304,105.5,-300.5</points>
<intersection>-304 1</intersection>
<intersection>-300.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-304,108.5,-304</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-300.5,105.5,-300.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-292,101,-286</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-286,101,-286</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-322.5,58.5,-237</points>
<intersection>-322.5 17</intersection>
<intersection>-311.5 15</intersection>
<intersection>-300 13</intersection>
<intersection>-289.5 11</intersection>
<intersection>-279 9</intersection>
<intersection>-267 7</intersection>
<intersection>-257 4</intersection>
<intersection>-246 5</intersection>
<intersection>-237 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-237,58.5,-237</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>55,-257,58.5,-257</points>
<connection>
<GID>9</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-246,58.5,-246</points>
<connection>
<GID>10</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54.5,-267,58.5,-267</points>
<connection>
<GID>8</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>55,-279,58.5,-279</points>
<connection>
<GID>89</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>55,-289.5,58.5,-289.5</points>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>55,-300,58.5,-300</points>
<connection>
<GID>5</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>55,-311.5,58.5,-311.5</points>
<connection>
<GID>6</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>55,-322.5,58.5,-322.5</points>
<connection>
<GID>7</GID>
<name>SEL_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-279,53.5,-240.5</points>
<connection>
<GID>10</GID>
<name>SEL_1</name></connection>
<connection>
<GID>8</GID>
<name>SEL_1</name></connection>
<intersection>-279 4</intersection>
<intersection>-257 2</intersection>
<intersection>-240.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-240.5,54,-240.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-257,54,-257</points>
<connection>
<GID>9</GID>
<name>SEL_1</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>53.5,-279,54,-279</points>
<connection>
<GID>89</GID>
<name>SEL_1</name></connection>
<intersection>53.5 0</intersection>
<intersection>54 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>54,-322.5,54,-279</points>
<connection>
<GID>7</GID>
<name>SEL_1</name></connection>
<connection>
<GID>6</GID>
<name>SEL_1</name></connection>
<connection>
<GID>5</GID>
<name>SEL_1</name></connection>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection>
<intersection>-279 4</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-305,83.5,-298</points>
<connection>
<GID>61</GID>
<name>load</name></connection>
<intersection>-298 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-298,83.5,-298</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-326.5,85.5,-316</points>
<connection>
<GID>61</GID>
<name>clear</name></connection>
<intersection>-326.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-326.5,85.5,-326.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-370,10.5,-361.5</points>
<connection>
<GID>62</GID>
<name>clear</name></connection>
<intersection>-370 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-370,10.5,-370</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-265.5,210,-258</points>
<intersection>-265.5 1</intersection>
<intersection>-258 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202,-265.5,210,-265.5</points>
<connection>
<GID>14</GID>
<name>ENABLE_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-258,210,-258</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-283,185.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_15</name></connection>
<intersection>-283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,-283,199,-283</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-286,186.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_14</name></connection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,-286,199,-286</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-290,187.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_13</name></connection>
<intersection>-290 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,-290,199,-290</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-294.5,188.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_12</name></connection>
<intersection>-294.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-294.5,199,-294.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-299,189.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_11</name></connection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,-299,199,-299</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-310.5,192.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_8</name></connection>
<intersection>-310.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,-310.5,198.5,-310.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175,-272.5,184,-272.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-271.5,179.5,-270.5</points>
<intersection>-271.5 1</intersection>
<intersection>-270.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-271.5,184,-271.5</points>
<connection>
<GID>14</GID>
<name>ADDRESS_1</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>175,-270.5,179.5,-270.5</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-270.5,179.5,-268.5</points>
<intersection>-270.5 1</intersection>
<intersection>-268.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-270.5,184,-270.5</points>
<connection>
<GID>14</GID>
<name>ADDRESS_2</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>175,-268.5,179.5,-268.5</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-269.5,179.5,-266.5</points>
<intersection>-269.5 1</intersection>
<intersection>-266.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-269.5,184,-269.5</points>
<connection>
<GID>14</GID>
<name>ADDRESS_3</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>175,-266.5,179.5,-266.5</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-328.5,29,-248.5</points>
<intersection>-328.5 2</intersection>
<intersection>-248.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-248.5,29,-248.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-328.5,51,-328.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-317.5,29,-246.5</points>
<intersection>-317.5 1</intersection>
<intersection>-246.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-317.5,51,-317.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-246.5,29,-246.5</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-306,29,-244.5</points>
<intersection>-306 1</intersection>
<intersection>-244.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-306,51,-306</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-244.5,29,-244.5</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-295.5,29,-242.5</points>
<intersection>-295.5 1</intersection>
<intersection>-242.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-295.5,51,-295.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-242.5,29,-242.5</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-285,29.5,-235</points>
<intersection>-285 1</intersection>
<intersection>-235 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-285,51,-285</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-235,29.5,-235</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-273,29,-233</points>
<intersection>-273 1</intersection>
<intersection>-233 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-273,50.5,-273</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-233,29,-233</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-263,29.5,-231</points>
<intersection>-263 1</intersection>
<intersection>-231 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-263,51,-263</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-231,29.5,-231</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-252,29,-229</points>
<intersection>-252 1</intersection>
<intersection>-229 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-252,50.5,-252</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-229,29,-229</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-303,191.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_9</name></connection>
<intersection>-303 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-303,199,-303</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-306.5,190.5,-276</points>
<connection>
<GID>14</GID>
<name>DATA_OUT_10</name></connection>
<intersection>-306.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,-306.5,199,-306.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>325.778,282.877,489.116,212.146</PageViewport></page 1>
<page 2>
<PageViewport>-129.882,41.9305,27.9978,-26.437</PageViewport></page 2>
<page 3>
<PageViewport>-138.149,45.3218,433.013,-202.012</PageViewport></page 3>
<page 4>
<PageViewport>77.4738,190.297,243.412,118.44</PageViewport></page 4>
<page 5>
<PageViewport>276.384,193.25,307.616,179.725</PageViewport></page 5>
<page 6>
<PageViewport>194.349,360.68,461.893,244.824</PageViewport></page 6>
<page 7>
<PageViewport>277.433,142.492,509.233,42.1143</PageViewport></page 7>
<page 8>
<PageViewport>84.8915,-47.6668,325.062,-151.669</PageViewport></page 8>
<page 9>
<PageViewport>597.038,118.247,768.872,43.8367</PageViewport></page 9></circuit>