<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-171.894,104.776,300.894,-144.913</PageViewport>
<gate>
<ID>2</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-17.5</position>
<input>
<ID>ENABLE_0</ID>20 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>55 </output>
<output>
<ID>OUT_1</ID>56 </output>
<output>
<ID>OUT_10</ID>65 </output>
<output>
<ID>OUT_11</ID>66 </output>
<output>
<ID>OUT_12</ID>67 </output>
<output>
<ID>OUT_13</ID>68 </output>
<output>
<ID>OUT_14</ID>69 </output>
<output>
<ID>OUT_15</ID>70 </output>
<output>
<ID>OUT_2</ID>57 </output>
<output>
<ID>OUT_3</ID>58 </output>
<output>
<ID>OUT_4</ID>59 </output>
<output>
<ID>OUT_5</ID>60 </output>
<output>
<ID>OUT_6</ID>61 </output>
<output>
<ID>OUT_7</ID>62 </output>
<output>
<ID>OUT_8</ID>63 </output>
<output>
<ID>OUT_9</ID>64 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>3</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>69,-40.5</position>
<input>
<ID>ENABLE_0</ID>19 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>12 </input>
<input>
<ID>IN_12</ID>13 </input>
<input>
<ID>IN_13</ID>14 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>16 </input>
<input>
<ID>IN_2</ID>3 </input>
<input>
<ID>IN_3</ID>4 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>6 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>8 </input>
<input>
<ID>IN_8</ID>9 </input>
<input>
<ID>IN_9</ID>10 </input>
<output>
<ID>OUT_0</ID>22 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_10</ID>44 </output>
<output>
<ID>OUT_11</ID>52 </output>
<output>
<ID>OUT_12</ID>45 </output>
<output>
<ID>OUT_13</ID>53 </output>
<output>
<ID>OUT_14</ID>46 </output>
<output>
<ID>OUT_15</ID>54 </output>
<output>
<ID>OUT_2</ID>40 </output>
<output>
<ID>OUT_3</ID>48 </output>
<output>
<ID>OUT_4</ID>41 </output>
<output>
<ID>OUT_5</ID>49 </output>
<output>
<ID>OUT_6</ID>42 </output>
<output>
<ID>OUT_7</ID>50 </output>
<output>
<ID>OUT_8</ID>43 </output>
<output>
<ID>OUT_9</ID>51 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>46.5,-4.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>16 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-35</position>
<output>
<ID>OUT_0</ID>9 </output>
<output>
<ID>OUT_1</ID>11 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>15 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>7</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-23</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>4 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>8 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>29,-47</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>7 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>1360</ID>
<type>AA_TOGGLE</type>
<position>20.5,118.5</position>
<output>
<ID>OUT_0</ID>1587 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>19.5,-36</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>19,-10</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>19,-22.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>19,-47.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BA_DECODER_2x4</type>
<position>60.5,-1</position>
<input>
<ID>ENABLE</ID>17 </input>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>55.5,0.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>51,-2.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>56,3.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>44.5,-2</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-36.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<input>
<ID>IN_2</ID>49 </input>
<input>
<ID>IN_3</ID>50 </input>
<input>
<ID>IN_B_0</ID>22 </input>
<input>
<ID>IN_B_1</ID>40 </input>
<input>
<ID>IN_B_2</ID>41 </input>
<input>
<ID>IN_B_3</ID>42 </input>
<output>
<ID>OUT_0</ID>71 </output>
<output>
<ID>OUT_1</ID>72 </output>
<output>
<ID>OUT_2</ID>73 </output>
<output>
<ID>OUT_3</ID>74 </output>
<output>
<ID>carry_out</ID>21 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_FULLADDER_4BIT</type>
<position>86.5,-52.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>53 </input>
<input>
<ID>IN_3</ID>54 </input>
<input>
<ID>IN_B_0</ID>43 </input>
<input>
<ID>IN_B_1</ID>44 </input>
<input>
<ID>IN_B_2</ID>45 </input>
<input>
<ID>IN_B_3</ID>46 </input>
<output>
<ID>OUT_0</ID>75 </output>
<output>
<ID>OUT_1</ID>76 </output>
<output>
<ID>OUT_2</ID>77 </output>
<output>
<ID>OUT_3</ID>78 </output>
<input>
<ID>carry_in</ID>21 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1186</ID>
<type>AA_LABEL</type>
<position>96.5,106</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>94,-29</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>94.5,-57.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1188</ID>
<type>AE_FULLADDER_4BIT</type>
<position>36.5,76</position>
<input>
<ID>IN_0</ID>1585 </input>
<input>
<ID>IN_1</ID>1587 </input>
<input>
<ID>IN_2</ID>1588 </input>
<input>
<ID>IN_3</ID>1589 </input>
<input>
<ID>IN_B_0</ID>1518 </input>
<input>
<ID>IN_B_1</ID>1529 </input>
<input>
<ID>IN_B_2</ID>1530 </input>
<input>
<ID>IN_B_3</ID>1531 </input>
<output>
<ID>OUT_0</ID>1591 </output>
<output>
<ID>OUT_1</ID>1592 </output>
<output>
<ID>OUT_2</ID>1593 </output>
<output>
<ID>OUT_3</ID>1663 </output>
<input>
<ID>carry_in</ID>1590 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1190</ID>
<type>AA_TOGGLE</type>
<position>-8,119</position>
<output>
<ID>OUT_0</ID>1589 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>80,-30</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>80.5,-36.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>80,-46</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>81,-53</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>82,-26</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1003</ID>
<type>AA_TOGGLE</type>
<position>32.5,119</position>
<output>
<ID>OUT_0</ID>1585 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>87,-22.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1390</ID>
<type>AA_TOGGLE</type>
<position>24.5,108</position>
<output>
<ID>OUT_0</ID>1529 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1004</ID>
<type>AA_TOGGLE</type>
<position>36.5,101.5</position>
<output>
<ID>OUT_0</ID>1518 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>82,-19</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>87,-15.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1392</ID>
<type>AA_LABEL</type>
<position>-2.5,123</position>
<gparam>LABEL_TEXT A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>82,-12</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>87,-8.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>82,-5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>87,-1.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_MUX_2x1</type>
<position>112,-13</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>94 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_MUX_2x1</type>
<position>112,-18</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>93 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1400</ID>
<type>AA_LABEL</type>
<position>0.5,105.5</position>
<gparam>LABEL_TEXT B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_MUX_2x1</type>
<position>112,-23</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>92 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1401</ID>
<type>AA_LABEL</type>
<position>7.5,122.5</position>
<gparam>LABEL_TEXT A6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_MUX_2x1</type>
<position>112,-28</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>91 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1402</ID>
<type>AA_LABEL</type>
<position>15.5,106</position>
<gparam>LABEL_TEXT B6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1209</ID>
<type>AA_TOGGLE</type>
<position>0.5,102</position>
<output>
<ID>OUT_0</ID>1531 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_MUX_2x1</type>
<position>112,-33</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>90 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1403</ID>
<type>AA_LABEL</type>
<position>26.5,123</position>
<gparam>LABEL_TEXT A5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_MUX_2x1</type>
<position>112,-38</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1404</ID>
<type>AA_LABEL</type>
<position>28.5,106</position>
<gparam>LABEL_TEXT B5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>112,-43</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>88 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1212</ID>
<type>AA_TOGGLE</type>
<position>7,118.5</position>
<output>
<ID>OUT_0</ID>1588 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_MUX_2x1</type>
<position>112,-48</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>87 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1407</ID>
<type>AE_FULLADDER_4BIT</type>
<position>63,75.5</position>
<input>
<ID>IN_0</ID>1512 </input>
<input>
<ID>IN_1</ID>1513 </input>
<input>
<ID>IN_2</ID>1514 </input>
<input>
<ID>IN_3</ID>1517 </input>
<input>
<ID>IN_B_0</ID>1466 </input>
<input>
<ID>IN_B_1</ID>1467 </input>
<input>
<ID>IN_B_2</ID>1468 </input>
<input>
<ID>IN_B_3</ID>1469 </input>
<output>
<ID>OUT_0</ID>1945 </output>
<output>
<ID>OUT_1</ID>1946 </output>
<output>
<ID>OUT_2</ID>1953 </output>
<output>
<ID>OUT_3</ID>1965 </output>
<output>
<ID>carry_out</ID>1590 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>134.5,-30</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>90 </input>
<input>
<ID>IN_4</ID>91 </input>
<input>
<ID>IN_5</ID>92 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>94 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1408</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>144.5,67.5</position>
<input>
<ID>IN_0</ID>1591 </input>
<input>
<ID>IN_1</ID>1592 </input>
<input>
<ID>IN_2</ID>1593 </input>
<input>
<ID>IN_3</ID>1663 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1024</ID>
<type>AA_TOGGLE</type>
<position>48,121</position>
<output>
<ID>OUT_0</ID>1517 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1027</ID>
<type>AA_TOGGLE</type>
<position>57.5,101.5</position>
<output>
<ID>OUT_0</ID>1469 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1031</ID>
<type>AA_TOGGLE</type>
<position>63.5,119</position>
<output>
<ID>OUT_0</ID>1514 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>112,-51.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1419</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>144.5,60.5</position>
<input>
<ID>IN_0</ID>1945 </input>
<input>
<ID>IN_1</ID>1946 </input>
<input>
<ID>IN_2</ID>1953 </input>
<input>
<ID>IN_3</ID>1965 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>113,-9</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1034</ID>
<type>AA_TOGGLE</type>
<position>71,101.5</position>
<output>
<ID>OUT_0</ID>1468 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1421</ID>
<type>AA_AND2</type>
<position>4.5,147.5</position>
<input>
<ID>IN_0</ID>1589 </input>
<input>
<ID>IN_1</ID>1531 </input>
<output>
<ID>OUT</ID>1966 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>126,-40</position>
<input>
<ID>N_in2</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1431</ID>
<type>AA_AND2</type>
<position>14.5,143.5</position>
<input>
<ID>IN_0</ID>1588 </input>
<input>
<ID>IN_1</ID>1530 </input>
<output>
<ID>OUT</ID>1967 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>128.5,-40</position>
<input>
<ID>N_in2</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1432</ID>
<type>AA_AND2</type>
<position>27.5,140</position>
<input>
<ID>IN_0</ID>1587 </input>
<input>
<ID>IN_1</ID>1529 </input>
<output>
<ID>OUT</ID>1975 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>131,-40</position>
<input>
<ID>N_in2</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1433</ID>
<type>AA_AND2</type>
<position>40.5,137.5</position>
<input>
<ID>IN_0</ID>1585 </input>
<input>
<ID>IN_1</ID>1518 </input>
<output>
<ID>OUT</ID>2004 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>133.5,-40</position>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1434</ID>
<type>AA_AND2</type>
<position>60,135</position>
<input>
<ID>IN_0</ID>1517 </input>
<input>
<ID>IN_1</ID>1469 </input>
<output>
<ID>OUT</ID>2005 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>136,-40</position>
<input>
<ID>N_in2</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>138.5,-40</position>
<input>
<ID>N_in2</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>141,-40</position>
<input>
<ID>N_in2</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1051</ID>
<type>AA_TOGGLE</type>
<position>75,119</position>
<output>
<ID>OUT_0</ID>1513 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>143.5,-40</position>
<input>
<ID>N_in2</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>143.5,-42</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>141,-42</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1441</ID>
<type>AA_AND2</type>
<position>72.5,132</position>
<input>
<ID>IN_0</ID>1514 </input>
<input>
<ID>IN_1</ID>1468 </input>
<output>
<ID>OUT</ID>2006 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>138.5,-42</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1442</ID>
<type>AA_AND2</type>
<position>86.5,129</position>
<input>
<ID>IN_0</ID>1513 </input>
<input>
<ID>IN_1</ID>1467 </input>
<output>
<ID>OUT</ID>2009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>136,-42</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1443</ID>
<type>AA_AND2</type>
<position>100,126</position>
<input>
<ID>IN_0</ID>1512 </input>
<input>
<ID>IN_1</ID>1466 </input>
<output>
<ID>OUT</ID>2010 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>133.5,-42</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1444</ID>
<type>AA_MUX_2x1</type>
<position>125,119.5</position>
<input>
<ID>IN_0</ID>1663 </input>
<input>
<ID>IN_1</ID>1966 </input>
<output>
<ID>OUT</ID>2051 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1445</ID>
<type>AA_MUX_2x1</type>
<position>125,114</position>
<input>
<ID>IN_0</ID>1593 </input>
<input>
<ID>IN_1</ID>1967 </input>
<output>
<ID>OUT</ID>2050 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>131,-42</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>128.5,-42</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1062</ID>
<type>AA_TOGGLE</type>
<position>83,101.5</position>
<output>
<ID>OUT_0</ID>1467 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>126,-42</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1064</ID>
<type>AA_TOGGLE</type>
<position>88.5,118.5</position>
<output>
<ID>OUT_0</ID>1512 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1066</ID>
<type>AA_TOGGLE</type>
<position>96,102</position>
<output>
<ID>OUT_0</ID>1466 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1456</ID>
<type>AA_MUX_2x1</type>
<position>125,109</position>
<input>
<ID>IN_0</ID>1592 </input>
<input>
<ID>IN_1</ID>1975 </input>
<output>
<ID>OUT</ID>2049 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1070</ID>
<type>AA_LABEL</type>
<position>40,123</position>
<gparam>LABEL_TEXT A4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1458</ID>
<type>AA_MUX_2x1</type>
<position>125,104</position>
<input>
<ID>IN_0</ID>1591 </input>
<input>
<ID>IN_1</ID>2004 </input>
<output>
<ID>OUT</ID>2048 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1459</ID>
<type>AA_MUX_2x1</type>
<position>125,99</position>
<input>
<ID>IN_0</ID>1965 </input>
<input>
<ID>IN_1</ID>2005 </input>
<output>
<ID>OUT</ID>2047 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1460</ID>
<type>AA_MUX_2x1</type>
<position>125,94</position>
<input>
<ID>IN_0</ID>1953 </input>
<input>
<ID>IN_1</ID>2006 </input>
<output>
<ID>OUT</ID>2013 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1461</ID>
<type>AA_MUX_2x1</type>
<position>125,89</position>
<input>
<ID>IN_0</ID>1946 </input>
<input>
<ID>IN_1</ID>2009 </input>
<output>
<ID>OUT</ID>2012 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1462</ID>
<type>AA_MUX_2x1</type>
<position>125,84</position>
<input>
<ID>IN_0</ID>1945 </input>
<input>
<ID>IN_1</ID>2010 </input>
<output>
<ID>OUT</ID>2011 </output>
<input>
<ID>SEL_0</ID>2061 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1463</ID>
<type>GA_LED</type>
<position>10,152</position>
<input>
<ID>N_in2</ID>1967 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1464</ID>
<type>GA_LED</type>
<position>-1.5,152</position>
<input>
<ID>N_in2</ID>1966 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1465</ID>
<type>GA_LED</type>
<position>20,151</position>
<input>
<ID>N_in2</ID>1975 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1079</ID>
<type>AA_LABEL</type>
<position>43,105.5</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1468</ID>
<type>GA_LED</type>
<position>32.5,150.5</position>
<input>
<ID>N_in2</ID>2004 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1470</ID>
<type>GA_LED</type>
<position>48.5,150</position>
<input>
<ID>N_in2</ID>2005 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1085</ID>
<type>AA_LABEL</type>
<position>55.5,122.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1472</ID>
<type>GA_LED</type>
<position>66,149</position>
<input>
<ID>N_in2</ID>2006 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1473</ID>
<type>GA_LED</type>
<position>79,149</position>
<input>
<ID>N_in2</ID>2009 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1087</ID>
<type>AA_LABEL</type>
<position>58,106</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1474</ID>
<type>GA_LED</type>
<position>103,148</position>
<input>
<ID>N_in2</ID>2010 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1475</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>143.5,101.5</position>
<input>
<ID>IN_0</ID>2011 </input>
<input>
<ID>IN_1</ID>2012 </input>
<input>
<ID>IN_2</ID>2013 </input>
<input>
<ID>IN_3</ID>2047 </input>
<input>
<ID>IN_4</ID>2048 </input>
<input>
<ID>IN_5</ID>2049 </input>
<input>
<ID>IN_6</ID>2050 </input>
<input>
<ID>IN_7</ID>2051 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1476</ID>
<type>AA_TOGGLE</type>
<position>121.5,123.5</position>
<output>
<ID>OUT_0</ID>2061 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1478</ID>
<type>AA_LABEL</type>
<position>57,183.5</position>
<gparam>LABEL_TEXT Original ALU</gparam>
<gparam>TEXT_HEIGHT 20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1480</ID>
<type>AA_LABEL</type>
<position>67.5,28.5</position>
<gparam>LABEL_TEXT Updated ALU</gparam>
<gparam>TEXT_HEIGHT 20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1294</ID>
<type>AA_TOGGLE</type>
<position>15,101.5</position>
<output>
<ID>OUT_0</ID>1530 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1120</ID>
<type>AA_LABEL</type>
<position>64.5,122.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1121</ID>
<type>AA_LABEL</type>
<position>71,106</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1149</ID>
<type>AA_LABEL</type>
<position>81,122.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1155</ID>
<type>AA_LABEL</type>
<position>83,105</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1156</ID>
<type>AA_LABEL</type>
<position>94.5,123</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-50,50.5,-48</points>
<intersection>-50 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-48,67,-48</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-50,50.5,-50</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-48,67,-25</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-47,50.5,-24</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection>
<intersection>-24 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-47,67,-47</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-26,50.5,-26</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-24,67,-24</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-48,50.5,-46</points>
<intersection>-48 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-46,67,-46</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-48,50.5,-48</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>67,-46,67,-23</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-45,50.5,-22</points>
<intersection>-45 1</intersection>
<intersection>-24 2</intersection>
<intersection>-22 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-45,67,-45</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-24,50.5,-24</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-22,67,-22</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-46,50.5,-44</points>
<intersection>-46 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-44,67,-44</points>
<connection>
<GID>3</GID>
<name>IN_4</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-46,50.5,-46</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-44,67,-21</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-43,50.5,-20</points>
<intersection>-43 1</intersection>
<intersection>-22 2</intersection>
<intersection>-20 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-43,67,-43</points>
<connection>
<GID>3</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-22,50.5,-22</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-20,67,-20</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-44,50.5,-42</points>
<intersection>-44 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-42,67,-42</points>
<connection>
<GID>3</GID>
<name>IN_6</name></connection>
<intersection>50.5 0</intersection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-44,50.5,-44</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-42,67,-19</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-41,50.5,-18</points>
<intersection>-41 1</intersection>
<intersection>-20 2</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-41,67,-41</points>
<connection>
<GID>3</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-20,50.5,-20</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-18,67,-18</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-40,50.5,-17</points>
<intersection>-40 1</intersection>
<intersection>-38 2</intersection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-40,67,-40</points>
<connection>
<GID>3</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-38,50.5,-38</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-17,67,-17</points>
<connection>
<GID>2</GID>
<name>IN_8</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-39,50.5,-14</points>
<intersection>-39 1</intersection>
<intersection>-16 4</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-39,67,-39</points>
<connection>
<GID>3</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-14,50.5,-14</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-16,67,-16</points>
<connection>
<GID>2</GID>
<name>IN_9</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-38,50.5,-15</points>
<intersection>-38 1</intersection>
<intersection>-36 2</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-38,67,-38</points>
<connection>
<GID>3</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-36,50.5,-36</points>
<connection>
<GID>6</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-15,67,-15</points>
<connection>
<GID>2</GID>
<name>IN_10</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-37,50.5,-12</points>
<intersection>-37 1</intersection>
<intersection>-14 3</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-37,67,-37</points>
<connection>
<GID>3</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-12,50.5,-12</points>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-14,67,-14</points>
<connection>
<GID>2</GID>
<name>IN_11</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-36,50.5,-13</points>
<intersection>-36 1</intersection>
<intersection>-34 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-36,67,-36</points>
<connection>
<GID>3</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-34,50.5,-34</points>
<connection>
<GID>6</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-13,67,-13</points>
<connection>
<GID>2</GID>
<name>IN_12</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-35,50.5,-10</points>
<intersection>-35 1</intersection>
<intersection>-12 3</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-35,67,-35</points>
<connection>
<GID>3</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-10,50.5,-10</points>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-12,67,-12</points>
<connection>
<GID>2</GID>
<name>IN_13</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1945</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,59.5,64.5,71.5</points>
<connection>
<GID>1407</GID>
<name>OUT_0</name></connection>
<intersection>59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,59.5,141.5,59.5</points>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection>
<intersection>123 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,59.5,123,83</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<intersection>59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-34,50.5,-11</points>
<intersection>-34 1</intersection>
<intersection>-32 2</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-34,67,-34</points>
<connection>
<GID>3</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-32,50.5,-32</points>
<connection>
<GID>6</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-11,67,-11</points>
<connection>
<GID>2</GID>
<name>IN_14</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,60.5,63.5,71.5</points>
<connection>
<GID>1407</GID>
<name>OUT_1</name></connection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,60.5,141.5,60.5</points>
<connection>
<GID>1419</GID>
<name>IN_1</name></connection>
<intersection>63.5 0</intersection>
<intersection>122 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>122,60.5,122,88</points>
<intersection>60.5 1</intersection>
<intersection>88 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,88,123,88</points>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection>
<intersection>122 2</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-33,50.5,-8</points>
<intersection>-33 1</intersection>
<intersection>-10 3</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-33,67,-33</points>
<connection>
<GID>3</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-8,50.5,-8</points>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-10,67,-10</points>
<connection>
<GID>2</GID>
<name>IN_15</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,0.5,57.5,0.5</points>
<connection>
<GID>15</GID>
<name>ENABLE</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,6,109,6</points>
<intersection>53 8</intersection>
<intersection>109 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>109,-45.5,109,6</points>
<intersection>-45.5 18</intersection>
<intersection>-40.5 19</intersection>
<intersection>-35.5 20</intersection>
<intersection>-30.5 21</intersection>
<intersection>-25.5 22</intersection>
<intersection>-20.5 23</intersection>
<intersection>-15.5 24</intersection>
<intersection>-10.5 25</intersection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>53,-2.5,53,6</points>
<intersection>-2.5 10</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>53,-2.5,57.5,-2.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>53 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>109,-45.5,112,-45.5</points>
<connection>
<GID>54</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>109,-40.5,112,-40.5</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>109,-35.5,112,-35.5</points>
<connection>
<GID>52</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>109,-30.5,112,-30.5</points>
<connection>
<GID>51</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>109,-25.5,112,-25.5</points>
<connection>
<GID>50</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>109,-20.5,112,-20.5</points>
<connection>
<GID>49</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>109,-15.5,112,-15.5</points>
<connection>
<GID>48</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>109,-10.5,112,-10.5</points>
<connection>
<GID>47</GID>
<name>SEL_0</name></connection>
<intersection>109 7</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-31.5,64.5,-2.5</points>
<intersection>-31.5 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-2.5,64.5,-2.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-31.5,69,-31.5</points>
<connection>
<GID>3</GID>
<name>ENABLE_0</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-8.5,69,-1.5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-1.5,69,-1.5</points>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-44.5,85.5,-44.5</points>
<connection>
<GID>25</GID>
<name>carry_out</name></connection>
<connection>
<GID>26</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-48,72.5,-31.5</points>
<intersection>-48 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-31.5,82.5,-31.5</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-48,72.5,-48</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,61.5,62.5,71.5</points>
<connection>
<GID>1407</GID>
<name>OUT_2</name></connection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,61.5,141.5,61.5</points>
<connection>
<GID>1419</GID>
<name>IN_2</name></connection>
<intersection>62.5 0</intersection>
<intersection>121 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>121,61.5,121,93</points>
<intersection>61.5 1</intersection>
<intersection>93 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>121,93,123,93</points>
<connection>
<GID>1460</GID>
<name>IN_0</name></connection>
<intersection>121 2</intersection></hsegment></shape></wire>
<wire>
<ID>1965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,62.5,61.5,71.5</points>
<connection>
<GID>1407</GID>
<name>OUT_3</name></connection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,62.5,141.5,62.5</points>
<connection>
<GID>1419</GID>
<name>IN_3</name></connection>
<intersection>61.5 0</intersection>
<intersection>120 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>120,62.5,120,98</points>
<intersection>62.5 1</intersection>
<intersection>98 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>120,98,123,98</points>
<connection>
<GID>1459</GID>
<name>IN_0</name></connection>
<intersection>120 2</intersection></hsegment></shape></wire>
<wire>
<ID>1966</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,147.5,-1.5,151</points>
<connection>
<GID>1464</GID>
<name>N_in2</name></connection>
<intersection>147.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,147.5,110,147.5</points>
<connection>
<GID>1421</GID>
<name>OUT</name></connection>
<intersection>-1.5 0</intersection>
<intersection>110 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>110,120.5,110,147.5</points>
<intersection>120.5 3</intersection>
<intersection>147.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>110,120.5,123,120.5</points>
<connection>
<GID>1444</GID>
<name>IN_1</name></connection>
<intersection>110 2</intersection></hsegment></shape></wire>
<wire>
<ID>1967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,143.5,10,151</points>
<connection>
<GID>1463</GID>
<name>N_in2</name></connection>
<intersection>143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,143.5,109,143.5</points>
<connection>
<GID>1431</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,115,109,143.5</points>
<intersection>115 4</intersection>
<intersection>143.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>109,115,123,115</points>
<connection>
<GID>1445</GID>
<name>IN_1</name></connection>
<intersection>109 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-46,73,-32.5</points>
<intersection>-46 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-32.5,82.5,-32.5</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-46,73,-46</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>1585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,80,34.5,138.5</points>
<connection>
<GID>1003</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1188</GID>
<name>IN_0</name></connection>
<intersection>138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,138.5,37.5,138.5</points>
<connection>
<GID>1433</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-44,73.5,-33.5</points>
<intersection>-44 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-33.5,82.5,-33.5</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-44,73.5,-44</points>
<connection>
<GID>3</GID>
<name>OUT_4</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-42,74,-34.5</points>
<intersection>-42 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-34.5,82.5,-34.5</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-42,74,-42</points>
<connection>
<GID>3</GID>
<name>OUT_6</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>1587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,80,33.5,86.5</points>
<connection>
<GID>1188</GID>
<name>IN_1</name></connection>
<intersection>86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,86.5,33.5,86.5</points>
<intersection>21.5 2</intersection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>21.5,86.5,21.5,141</points>
<intersection>86.5 1</intersection>
<intersection>118.5 5</intersection>
<intersection>141 7</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>21.5,118.5,22.5,118.5</points>
<connection>
<GID>1360</GID>
<name>OUT_0</name></connection>
<intersection>21.5 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,141,24.5,141</points>
<connection>
<GID>1432</GID>
<name>IN_0</name></connection>
<intersection>21.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-47.5,76,-40</points>
<intersection>-47.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-47.5,82.5,-47.5</points>
<connection>
<GID>26</GID>
<name>IN_B_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-40,76,-40</points>
<connection>
<GID>3</GID>
<name>OUT_8</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>1588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,80,32.5,88.5</points>
<connection>
<GID>1188</GID>
<name>IN_2</name></connection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,88.5,32.5,88.5</points>
<intersection>12 2</intersection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>12,88.5,12,119</points>
<intersection>88.5 1</intersection>
<intersection>119 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>9,119,12,119</points>
<intersection>9 6</intersection>
<intersection>9.5 7</intersection>
<intersection>12 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>9,118.5,9,119</points>
<connection>
<GID>1212</GID>
<name>OUT_0</name></connection>
<intersection>119 5</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>9.5,119,9.5,144.5</points>
<intersection>119 5</intersection>
<intersection>144.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>9.5,144.5,11.5,144.5</points>
<connection>
<GID>1431</GID>
<name>IN_0</name></connection>
<intersection>9.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-48.5,75.5,-38</points>
<intersection>-48.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-48.5,82.5,-48.5</points>
<connection>
<GID>26</GID>
<name>IN_B_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-38,75.5,-38</points>
<connection>
<GID>3</GID>
<name>OUT_10</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,140,20,150</points>
<connection>
<GID>1465</GID>
<name>N_in2</name></connection>
<intersection>140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,140,108,140</points>
<connection>
<GID>1432</GID>
<name>OUT</name></connection>
<intersection>20 0</intersection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,110,108,140</points>
<intersection>110 3</intersection>
<intersection>140 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>108,110,123,110</points>
<connection>
<GID>1456</GID>
<name>IN_1</name></connection>
<intersection>108 2</intersection></hsegment></shape></wire>
<wire>
<ID>1589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,80,31.5,86</points>
<connection>
<GID>1188</GID>
<name>IN_3</name></connection>
<intersection>86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,86,31.5,86</points>
<intersection>-4 2</intersection>
<intersection>31.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-4,86,-4,115.5</points>
<intersection>86 1</intersection>
<intersection>115.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,115.5,0,115.5</points>
<intersection>-4 2</intersection>
<intersection>0 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>0,115.5,0,148.5</points>
<intersection>115.5 3</intersection>
<intersection>119 6</intersection>
<intersection>148.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>0,148.5,1.5,148.5</points>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection>
<intersection>0 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6,119,0,119</points>
<connection>
<GID>1190</GID>
<name>OUT_0</name></connection>
<intersection>0 4</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-49.5,75,-36</points>
<intersection>-49.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-49.5,82.5,-49.5</points>
<connection>
<GID>26</GID>
<name>IN_B_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-36,75,-36</points>
<connection>
<GID>3</GID>
<name>OUT_12</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>1590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,76.5,55,76.5</points>
<connection>
<GID>1407</GID>
<name>carry_out</name></connection>
<intersection>44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,76.5,44.5,77</points>
<connection>
<GID>1188</GID>
<name>carry_in</name></connection>
<intersection>76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-50.5,74.5,-34</points>
<intersection>-50.5 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-50.5,82.5,-50.5</points>
<connection>
<GID>26</GID>
<name>IN_B_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-34,74.5,-34</points>
<connection>
<GID>3</GID>
<name>OUT_14</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,66.5,38,72</points>
<connection>
<GID>1188</GID>
<name>OUT_0</name></connection>
<intersection>66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,66.5,141.5,66.5</points>
<connection>
<GID>1408</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection>
<intersection>119 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119,66.5,119,103</points>
<intersection>66.5 1</intersection>
<intersection>103 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119,103,123,103</points>
<connection>
<GID>1458</GID>
<name>IN_0</name></connection>
<intersection>119 2</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-47,76.5,-38.5</points>
<intersection>-47 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-38.5,82.5,-38.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-47,76.5,-47</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,67.5,37,72</points>
<connection>
<GID>1188</GID>
<name>OUT_1</name></connection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,67.5,141.5,67.5</points>
<connection>
<GID>1408</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection>
<intersection>118 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>118,67.5,118,108</points>
<intersection>67.5 1</intersection>
<intersection>108 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>118,108,123,108</points>
<connection>
<GID>1456</GID>
<name>IN_0</name></connection>
<intersection>118 2</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-45,76.5,-39.5</points>
<intersection>-45 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-39.5,82.5,-39.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-45,76.5,-45</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,68.5,36,72</points>
<connection>
<GID>1188</GID>
<name>OUT_2</name></connection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,68.5,141.5,68.5</points>
<connection>
<GID>1408</GID>
<name>IN_2</name></connection>
<intersection>36 0</intersection>
<intersection>117 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>117,68.5,117,113</points>
<intersection>68.5 1</intersection>
<intersection>113 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>117,113,123,113</points>
<connection>
<GID>1445</GID>
<name>IN_0</name></connection>
<intersection>117 2</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-43,76.5,-40.5</points>
<intersection>-43 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-40.5,82.5,-40.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-43,76.5,-43</points>
<connection>
<GID>3</GID>
<name>OUT_5</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-41.5,76.5,-41</points>
<intersection>-41.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-41.5,82.5,-41.5</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-41,76.5,-41</points>
<connection>
<GID>3</GID>
<name>OUT_7</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-54.5,78.5,-39</points>
<intersection>-54.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-54.5,82.5,-54.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-39,78.5,-39</points>
<connection>
<GID>3</GID>
<name>OUT_9</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-55.5,78,-37</points>
<intersection>-55.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-55.5,82.5,-55.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-37,78,-37</points>
<connection>
<GID>3</GID>
<name>OUT_11</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-56.5,77.5,-35</points>
<intersection>-56.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-56.5,82.5,-56.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-35,77.5,-35</points>
<connection>
<GID>3</GID>
<name>OUT_13</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-57.5,77,-33</points>
<intersection>-57.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-57.5,82.5,-57.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-33,77,-33</points>
<connection>
<GID>3</GID>
<name>OUT_15</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-27,72,-25</points>
<intersection>-27 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-27,79,-27</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-25,72,-25</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-25,79,-25</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-25,71,-24</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-23.5,74.5,-23</points>
<intersection>-23.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-23.5,84,-23.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-23,74.5,-23</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-21.5,84,-21.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-22,71,-21.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-20,79,-20</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-21,71,-20</points>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-20,72,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-18,79,-18</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-20,72,-20</points>
<connection>
<GID>2</GID>
<name>OUT_5</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-19,73,-16.5</points>
<intersection>-19 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-16.5,84,-16.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-19,73,-19</points>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-18,72.5,-14.5</points>
<intersection>-18 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-14.5,84,-14.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-18,72.5,-18</points>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-17,72,-13</points>
<intersection>-17 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-13,79,-13</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-17,72,-17</points>
<connection>
<GID>2</GID>
<name>OUT_8</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-16,72,-11</points>
<intersection>-16 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-11,79,-11</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-16,72,-16</points>
<connection>
<GID>2</GID>
<name>OUT_9</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-15,72.5,-9.5</points>
<intersection>-15 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-9.5,84,-9.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-15,72.5,-15</points>
<connection>
<GID>2</GID>
<name>OUT_10</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-14,72.5,-7.5</points>
<intersection>-14 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-7.5,84,-7.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-14,72.5,-14</points>
<connection>
<GID>2</GID>
<name>OUT_11</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-13,72,-6</points>
<intersection>-13 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-6,79,-6</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-13,72,-13</points>
<connection>
<GID>2</GID>
<name>OUT_12</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-12,72,-4</points>
<intersection>-12 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-4,79,-4</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-12,72,-12</points>
<connection>
<GID>2</GID>
<name>OUT_13</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-11,71.5,-2.5</points>
<intersection>-11 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-2.5,84,-2.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-11,71.5,-11</points>
<connection>
<GID>2</GID>
<name>OUT_14</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-10,71,-0.5</points>
<connection>
<GID>2</GID>
<name>OUT_15</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-0.5,84,-0.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-49,100,-35</points>
<intersection>-49 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-49,110,-49</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-35,100,-35</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-44,100,-36</points>
<intersection>-44 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-44,110,-44</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-36,100,-36</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-39,100,-37</points>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-39,110,-39</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-37,100,-37</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,137.5,32.5,149.5</points>
<connection>
<GID>1468</GID>
<name>N_in2</name></connection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,137.5,107,137.5</points>
<connection>
<GID>1433</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection>
<intersection>107 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>107,105,107,137.5</points>
<intersection>105 3</intersection>
<intersection>137.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,105,123,105</points>
<connection>
<GID>1458</GID>
<name>IN_1</name></connection>
<intersection>107 2</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-38,100,-34</points>
<intersection>-38 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-34,110,-34</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-38,100,-38</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,135,48.5,149</points>
<connection>
<GID>1470</GID>
<name>N_in2</name></connection>
<intersection>135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,135,106,135</points>
<connection>
<GID>1434</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection>
<intersection>106 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>106,100,106,135</points>
<intersection>100 3</intersection>
<intersection>135 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>106,100,123,100</points>
<connection>
<GID>1459</GID>
<name>IN_1</name></connection>
<intersection>106 2</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-51,100,-29</points>
<intersection>-51 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-29,110,-29</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-51,100,-51</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,132,66,148</points>
<connection>
<GID>1472</GID>
<name>N_in2</name></connection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,132,105,132</points>
<connection>
<GID>1441</GID>
<name>OUT</name></connection>
<intersection>66 0</intersection>
<intersection>105 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>105,95,105,132</points>
<intersection>95 3</intersection>
<intersection>132 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>105,95,123,95</points>
<connection>
<GID>1460</GID>
<name>IN_1</name></connection>
<intersection>105 2</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-52,100,-24</points>
<intersection>-52 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-24,110,-24</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-52,100,-52</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-53,100,-19</points>
<intersection>-53 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-19,110,-19</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-53,100,-53</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-54,100,-14</points>
<intersection>-54 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-14,110,-14</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-54,100,-54</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,129,79,148</points>
<connection>
<GID>1473</GID>
<name>N_in2</name></connection>
<intersection>129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,129,104,129</points>
<connection>
<GID>1442</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection>
<intersection>104 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>104,90,104,129</points>
<intersection>90 3</intersection>
<intersection>129 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>104,90,123,90</points>
<connection>
<GID>1461</GID>
<name>IN_1</name></connection>
<intersection>104 2</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-47,97.5,-26</points>
<intersection>-47 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-47,110,-47</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-26,97.5,-26</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,85,103,147</points>
<connection>
<GID>1443</GID>
<name>OUT</name></connection>
<connection>
<GID>1474</GID>
<name>N_in2</name></connection>
<intersection>85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,85,123,85</points>
<connection>
<GID>1462</GID>
<name>IN_1</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-42,100,-22.5</points>
<intersection>-42 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-22.5,100,-22.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-42,110,-42</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,84,132.5,98.5</points>
<intersection>84 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,98.5,138.5,98.5</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,84,132.5,84</points>
<connection>
<GID>1462</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-37,97.5,-19</points>
<intersection>-37 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-19,97.5,-19</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-37,110,-37</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,89,132.5,99.5</points>
<intersection>89 2</intersection>
<intersection>99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,99.5,138.5,99.5</points>
<connection>
<GID>1475</GID>
<name>IN_1</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,89,132.5,89</points>
<connection>
<GID>1461</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-32,100,-15.5</points>
<intersection>-32 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-15.5,100,-15.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-32,110,-32</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>2013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,94,132.5,100.5</points>
<intersection>94 2</intersection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,100.5,138.5,100.5</points>
<connection>
<GID>1475</GID>
<name>IN_2</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,94,132.5,94</points>
<connection>
<GID>1460</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-27,97.5,-12</points>
<intersection>-27 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-12,97.5,-12</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-27,110,-27</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-22,100,-8.5</points>
<intersection>-22 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-8.5,100,-8.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-22,110,-22</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-17,97.5,-5</points>
<intersection>-17 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-5,97.5,-5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-17,110,-17</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-12,100,-1.5</points>
<intersection>-12 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-1.5,100,-1.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-12,110,-12</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-48,121.5,-33</points>
<intersection>-48 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-33,129.5,-33</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection>
<intersection>122.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-48,121.5,-48</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>122.5,-38.5,122.5,-33</points>
<intersection>-38.5 8</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>122.5,-38.5,143.5,-38.5</points>
<intersection>122.5 7</intersection>
<intersection>143.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>143.5,-39,143.5,-38.5</points>
<connection>
<GID>86</GID>
<name>N_in2</name></connection>
<intersection>-38.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-43,121.5,-32</points>
<intersection>-43 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-32,129.5,-32</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection>
<intersection>123 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-43,121.5,-43</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123,-38,123,-32</points>
<intersection>-38 8</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123,-38,141,-38</points>
<intersection>123 7</intersection>
<intersection>141 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>141,-39,141,-38</points>
<connection>
<GID>85</GID>
<name>N_in2</name></connection>
<intersection>-38 8</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-38,121.5,-31</points>
<intersection>-38 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-31,129.5,-31</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>121.5 0</intersection>
<intersection>123.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-38,121.5,-38</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>123.5,-37.5,123.5,-31</points>
<intersection>-37.5 8</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>123.5,-37.5,138.5,-37.5</points>
<intersection>123.5 7</intersection>
<intersection>138.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>138.5,-39,138.5,-37.5</points>
<connection>
<GID>84</GID>
<name>N_in2</name></connection>
<intersection>-37.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-33,121.5,-30</points>
<intersection>-33 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-30,129.5,-30</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>121.5 0</intersection>
<intersection>124 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-33,121.5,-33</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124,-37,124,-30</points>
<intersection>-37 9</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124,-37,136,-37</points>
<intersection>124 8</intersection>
<intersection>136 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>136,-39,136,-37</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>-37 9</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-29,121.5,-28</points>
<intersection>-29 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-29,129.5,-29</points>
<connection>
<GID>56</GID>
<name>IN_4</name></connection>
<intersection>121.5 0</intersection>
<intersection>124.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-28,121.5,-28</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>124.5,-36.5,124.5,-29</points>
<intersection>-36.5 9</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>124.5,-36.5,133.5,-36.5</points>
<intersection>124.5 8</intersection>
<intersection>133.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>133.5,-39,133.5,-36.5</points>
<connection>
<GID>82</GID>
<name>N_in2</name></connection>
<intersection>-36.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-28,121.5,-23</points>
<intersection>-28 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-28,129.5,-28</points>
<connection>
<GID>56</GID>
<name>IN_5</name></connection>
<intersection>121.5 0</intersection>
<intersection>125 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-23,121.5,-23</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125,-36,125,-28</points>
<intersection>-36 8</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125,-36,131,-36</points>
<intersection>125 7</intersection>
<intersection>131 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>131,-39,131,-36</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<intersection>-36 8</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-27,121.5,-18</points>
<intersection>-27 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-27,129.5,-27</points>
<connection>
<GID>56</GID>
<name>IN_6</name></connection>
<intersection>121.5 0</intersection>
<intersection>125.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114,-18,121.5,-18</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>125.5,-35.5,125.5,-27</points>
<intersection>-35.5 8</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>125.5,-35.5,128.5,-35.5</points>
<intersection>125.5 7</intersection>
<intersection>128.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>128.5,-39,128.5,-35.5</points>
<connection>
<GID>80</GID>
<name>N_in2</name></connection>
<intersection>-35.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-26,121.5,-13</points>
<intersection>-26 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114,-13,121.5,-13</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-26,129.5,-26</points>
<connection>
<GID>56</GID>
<name>IN_7</name></connection>
<intersection>121.5 0</intersection>
<intersection>126 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>126,-39,126,-26</points>
<connection>
<GID>79</GID>
<name>N_in2</name></connection>
<intersection>-26 2</intersection></vsegment></shape></wire>
<wire>
<ID>1466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,80,97,80</points>
<intersection>68 4</intersection>
<intersection>97 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>97,80,97,125</points>
<connection>
<GID>1443</GID>
<name>IN_1</name></connection>
<intersection>80 1</intersection>
<intersection>102 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>68,79.5,68,80</points>
<connection>
<GID>1407</GID>
<name>IN_B_0</name></connection>
<intersection>80 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>97,102,98,102</points>
<connection>
<GID>1066</GID>
<name>OUT_0</name></connection>
<intersection>97 2</intersection></hsegment></shape></wire>
<wire>
<ID>1467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,79.5,67,83</points>
<connection>
<GID>1407</GID>
<name>IN_B_1</name></connection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,83,83.5,83</points>
<intersection>67 0</intersection>
<intersection>83.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,83,83.5,128</points>
<connection>
<GID>1442</GID>
<name>IN_1</name></connection>
<intersection>83 1</intersection>
<intersection>101.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>83.5,101.5,85,101.5</points>
<connection>
<GID>1062</GID>
<name>OUT_0</name></connection>
<intersection>83.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2047</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,99,132.5,101.5</points>
<intersection>99 2</intersection>
<intersection>101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,101.5,138.5,101.5</points>
<connection>
<GID>1475</GID>
<name>IN_3</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,99,132.5,99</points>
<connection>
<GID>1459</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,79.5,66,84</points>
<connection>
<GID>1407</GID>
<name>IN_B_2</name></connection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,84,69.5,84</points>
<intersection>66 0</intersection>
<intersection>69.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>69.5,84,69.5,131</points>
<connection>
<GID>1441</GID>
<name>IN_1</name></connection>
<intersection>84 1</intersection>
<intersection>101.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>69.5,101.5,73,101.5</points>
<connection>
<GID>1034</GID>
<name>OUT_0</name></connection>
<intersection>69.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2048</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,102.5,132.5,104</points>
<intersection>102.5 1</intersection>
<intersection>104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,102.5,138.5,102.5</points>
<connection>
<GID>1475</GID>
<name>IN_4</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,104,132.5,104</points>
<connection>
<GID>1458</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,79.5,65,83.5</points>
<connection>
<GID>1407</GID>
<name>IN_B_3</name></connection>
<intersection>83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,83.5,65,83.5</points>
<intersection>59.5 2</intersection>
<intersection>65 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>59.5,83.5,59.5,134</points>
<connection>
<GID>1027</GID>
<name>OUT_0</name></connection>
<intersection>83.5 1</intersection>
<intersection>134 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,134,59.5,134</points>
<connection>
<GID>1434</GID>
<name>IN_1</name></connection>
<intersection>59.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,103.5,132.5,109</points>
<intersection>103.5 1</intersection>
<intersection>109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,103.5,138.5,103.5</points>
<connection>
<GID>1475</GID>
<name>IN_5</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,109,132.5,109</points>
<connection>
<GID>1456</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,69.5,35,72</points>
<connection>
<GID>1188</GID>
<name>OUT_3</name></connection>
<intersection>69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,69.5,141.5,69.5</points>
<connection>
<GID>1408</GID>
<name>IN_3</name></connection>
<intersection>35 0</intersection>
<intersection>116 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>116,69.5,116,118.5</points>
<intersection>69.5 1</intersection>
<intersection>118.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>116,118.5,123,118.5</points>
<connection>
<GID>1444</GID>
<name>IN_0</name></connection>
<intersection>116 2</intersection></hsegment></shape></wire>
<wire>
<ID>2050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,104.5,132.5,114</points>
<intersection>104.5 1</intersection>
<intersection>114 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,104.5,138.5,104.5</points>
<connection>
<GID>1475</GID>
<name>IN_6</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,114,132.5,114</points>
<connection>
<GID>1445</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,105.5,132.5,119.5</points>
<intersection>105.5 1</intersection>
<intersection>119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,105.5,138.5,105.5</points>
<connection>
<GID>1475</GID>
<name>IN_7</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,119.5,132.5,119.5</points>
<connection>
<GID>1444</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2061</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,86.5,125,123.5</points>
<connection>
<GID>1462</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1461</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1460</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1459</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1458</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1456</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1445</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1444</GID>
<name>SEL_0</name></connection>
<intersection>123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,123.5,125,123.5</points>
<connection>
<GID>1476</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>1512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,79.5,61,86.5</points>
<connection>
<GID>1407</GID>
<name>IN_0</name></connection>
<intersection>86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,86.5,93,86.5</points>
<intersection>61 0</intersection>
<intersection>93 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>93,86.5,93,127</points>
<intersection>86.5 1</intersection>
<intersection>118.5 5</intersection>
<intersection>127 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>90.5,118.5,93,118.5</points>
<connection>
<GID>1064</GID>
<name>OUT_0</name></connection>
<intersection>93 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>93,127,97,127</points>
<connection>
<GID>1443</GID>
<name>IN_0</name></connection>
<intersection>93 2</intersection></hsegment></shape></wire>
<wire>
<ID>1513</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,79.5,60,88</points>
<connection>
<GID>1407</GID>
<name>IN_1</name></connection>
<intersection>88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,88,78.5,88</points>
<intersection>60 0</intersection>
<intersection>78.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>78.5,88,78.5,130</points>
<intersection>88 1</intersection>
<intersection>119 5</intersection>
<intersection>130 7</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>77,119,78.5,119</points>
<connection>
<GID>1051</GID>
<name>OUT_0</name></connection>
<intersection>78.5 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>78.5,130,83.5,130</points>
<connection>
<GID>1442</GID>
<name>IN_0</name></connection>
<intersection>78.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1514</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,79.5,59,89.5</points>
<connection>
<GID>1407</GID>
<name>IN_2</name></connection>
<intersection>89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,89.5,68,89.5</points>
<intersection>59 0</intersection>
<intersection>68 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>68,89.5,68,133</points>
<intersection>89.5 1</intersection>
<intersection>119 3</intersection>
<intersection>133 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>65.5,119,68,119</points>
<connection>
<GID>1031</GID>
<name>OUT_0</name></connection>
<intersection>68 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>68,133,69.5,133</points>
<connection>
<GID>1441</GID>
<name>IN_0</name></connection>
<intersection>68 2</intersection></hsegment></shape></wire>
<wire>
<ID>1517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,79.5,58,84.5</points>
<connection>
<GID>1407</GID>
<name>IN_3</name></connection>
<intersection>84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,84.5,58,84.5</points>
<intersection>54.5 2</intersection>
<intersection>58 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>54.5,84.5,54.5,115.5</points>
<intersection>84.5 1</intersection>
<intersection>115.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>50,115.5,54.5,115.5</points>
<intersection>50 4</intersection>
<intersection>54.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,115.5,50,136</points>
<connection>
<GID>1024</GID>
<name>OUT_0</name></connection>
<intersection>115.5 3</intersection>
<intersection>136 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50,136,57,136</points>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection>
<intersection>50 4</intersection></hsegment></shape></wire>
<wire>
<ID>1518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,80,46.5,100</points>
<intersection>80 2</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,100,46.5,100</points>
<intersection>38.5 3</intersection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,80,46.5,80</points>
<connection>
<GID>1188</GID>
<name>IN_B_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38.5,100,38.5,136.5</points>
<connection>
<GID>1004</GID>
<name>OUT_0</name></connection>
<intersection>100 1</intersection>
<intersection>136.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,136.5,38.5,136.5</points>
<connection>
<GID>1433</GID>
<name>IN_1</name></connection>
<intersection>38.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,80,40.5,82</points>
<connection>
<GID>1188</GID>
<name>IN_B_1</name></connection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,82,40.5,82</points>
<intersection>30.5 2</intersection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>30.5,82,30.5,108</points>
<intersection>82 1</intersection>
<intersection>108 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,108,30.5,108</points>
<connection>
<GID>1390</GID>
<name>OUT_0</name></connection>
<intersection>26.5 4</intersection>
<intersection>30.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26.5,108,26.5,139</points>
<intersection>108 3</intersection>
<intersection>139 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>24.5,139,26.5,139</points>
<connection>
<GID>1432</GID>
<name>IN_1</name></connection>
<intersection>26.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,80,39.5,85.5</points>
<connection>
<GID>1188</GID>
<name>IN_B_2</name></connection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,85.5,39.5,85.5</points>
<intersection>17 2</intersection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>17,85.5,17,142.5</points>
<connection>
<GID>1294</GID>
<name>OUT_0</name></connection>
<intersection>85.5 1</intersection>
<intersection>142.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>11.5,142.5,17,142.5</points>
<connection>
<GID>1431</GID>
<name>IN_1</name></connection>
<intersection>17 2</intersection></hsegment></shape></wire>
<wire>
<ID>1531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,80,38.5,83</points>
<connection>
<GID>1188</GID>
<name>IN_B_3</name></connection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,83,38.5,83</points>
<intersection>2.5 2</intersection>
<intersection>38.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>2.5,83,2.5,146.5</points>
<connection>
<GID>1209</GID>
<name>OUT_0</name></connection>
<intersection>83 1</intersection>
<intersection>146.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1.5,146.5,2.5,146.5</points>
<connection>
<GID>1421</GID>
<name>IN_1</name></connection>
<intersection>2.5 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-21.771,-24.7071,214.521,-149.498</PageViewport>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>166.5,-34</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>166.5,-45</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AE_REGISTER8</type>
<position>109.5,-45</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>128 </output>
<output>
<ID>OUT_1</ID>127 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>125 </output>
<output>
<ID>OUT_4</ID>124 </output>
<output>
<ID>OUT_5</ID>123 </output>
<output>
<ID>OUT_6</ID>122 </output>
<output>
<ID>OUT_7</ID>121 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>168 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_REGISTER8</type>
<position>109.5,-58</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>144 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>133 </output>
<output>
<ID>OUT_4</ID>132 </output>
<output>
<ID>OUT_5</ID>131 </output>
<output>
<ID>OUT_6</ID>130 </output>
<output>
<ID>OUT_7</ID>129 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>169 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>60</ID>
<type>AE_MUX_4x1</type>
<position>135,-7.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>136 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>AE_MUX_4x1</type>
<position>135,-18.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>122 </input>
<input>
<ID>IN_2</ID>114 </input>
<input>
<ID>IN_3</ID>106 </input>
<output>
<ID>OUT</ID>137 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_MUX_4x1</type>
<position>135,-29.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT</ID>138 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_MUX_4x1</type>
<position>135,-39</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>108 </input>
<output>
<ID>OUT</ID>139 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_MUX_4x1</type>
<position>135,-50</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>117 </input>
<input>
<ID>IN_3</ID>109 </input>
<output>
<ID>OUT</ID>140 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_MUX_4x1</type>
<position>135,-61</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_MUX_4x1</type>
<position>135,-71.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>119 </input>
<input>
<ID>IN_3</ID>111 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_MUX_4x1</type>
<position>135,-82.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>112 </input>
<output>
<ID>OUT</ID>143 </output>
<input>
<ID>SEL_0</ID>146 </input>
<input>
<ID>SEL_1</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>70</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>167,-40</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>140 </input>
<input>
<ID>IN_4</ID>139 </input>
<input>
<ID>IN_5</ID>138 </input>
<input>
<ID>IN_6</ID>137 </input>
<input>
<ID>IN_7</ID>136 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>71</ID>
<type>DD_KEYPAD_HEX</type>
<position>76.5,-22.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<output>
<ID>OUT_1</ID>147 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>BB_CLOCK</type>
<position>98,-66.5</position>
<output>
<ID>CLK</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>110.5,-11.5</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>110.5,-24.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>110.5,-38</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>110.5,-51</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>75,-15.5</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>DD_KEYPAD_HEX</type>
<position>76.5,-36.5</position>
<output>
<ID>OUT_0</ID>156 </output>
<output>
<ID>OUT_1</ID>157 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-7.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>148 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-18.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>122 </input>
<input>
<ID>IN_2</ID>114 </input>
<input>
<ID>IN_3</ID>106 </input>
<output>
<ID>OUT</ID>149 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-29.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>123 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>107 </input>
<output>
<ID>OUT</ID>150 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-39</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>116 </input>
<input>
<ID>IN_3</ID>108 </input>
<output>
<ID>OUT</ID>151 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-50</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>125 </input>
<input>
<ID>IN_2</ID>117 </input>
<input>
<ID>IN_3</ID>109 </input>
<output>
<ID>OUT</ID>152 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-61</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT</ID>153 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-71.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>119 </input>
<input>
<ID>IN_3</ID>111 </input>
<output>
<ID>OUT</ID>154 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_MUX_4x1</type>
<position>147.5,-82.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>112 </input>
<output>
<ID>OUT</ID>155 </output>
<input>
<ID>SEL_0</ID>156 </input>
<input>
<ID>SEL_1</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>103</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>167,-51</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<input>
<ID>IN_4</ID>151 </input>
<input>
<ID>IN_5</ID>150 </input>
<input>
<ID>IN_6</ID>149 </input>
<input>
<ID>IN_7</ID>148 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>75,-29.5</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>DD_KEYPAD_HEX</type>
<position>92.5,-36</position>
<output>
<ID>OUT_0</ID>161 </output>
<output>
<ID>OUT_1</ID>160 </output>
<output>
<ID>OUT_2</ID>159 </output>
<output>
<ID>OUT_3</ID>158 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>106</ID>
<type>DD_KEYPAD_HEX</type>
<position>92.5,-48</position>
<output>
<ID>OUT_0</ID>165 </output>
<output>
<ID>OUT_1</ID>164 </output>
<output>
<ID>OUT_2</ID>163 </output>
<output>
<ID>OUT_3</ID>162 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>92.5,-29</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>BA_DECODER_2x4</type>
<position>94.5,-3</position>
<input>
<ID>ENABLE</ID>170 </input>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT_0</ID>166 </output>
<output>
<ID>OUT_1</ID>167 </output>
<output>
<ID>OUT_2</ID>168 </output>
<output>
<ID>OUT_3</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>88.5,-2.5</position>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>86,-1</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>DD_KEYPAD_HEX</type>
<position>89.5,-15.5</position>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>172 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>90,-8.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AE_REGISTER8</type>
<position>109.5,-18.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>112 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>110 </output>
<output>
<ID>OUT_3</ID>109 </output>
<output>
<ID>OUT_4</ID>108 </output>
<output>
<ID>OUT_5</ID>107 </output>
<output>
<ID>OUT_6</ID>106 </output>
<output>
<ID>OUT_7</ID>105 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>166 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_REGISTER8</type>
<position>109.5,-31.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>161 </input>
<input>
<ID>IN_5</ID>160 </input>
<input>
<ID>IN_6</ID>159 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT_0</ID>120 </output>
<output>
<ID>OUT_1</ID>119 </output>
<output>
<ID>OUT_2</ID>118 </output>
<output>
<ID>OUT_3</ID>117 </output>
<output>
<ID>OUT_4</ID>116 </output>
<output>
<ID>OUT_5</ID>115 </output>
<output>
<ID>OUT_6</ID>114 </output>
<output>
<ID>OUT_7</ID>113 </output>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>load</ID>167 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>120,6</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-14.5,131.5,-14.5</points>
<connection>
<GID>113</GID>
<name>OUT_7</name></connection>
<intersection>131.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131.5,-14.5,131.5,-4.5</points>
<intersection>-14.5 1</intersection>
<intersection>-4.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>131.5,-4.5,144.5,-4.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<intersection>131.5 4</intersection>
<intersection>143 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>143,-10.5,143,-4.5</points>
<intersection>-10.5 8</intersection>
<intersection>-4.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>143,-10.5,144.5,-10.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>143 6</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-15.5,144.5,-15.5</points>
<connection>
<GID>113</GID>
<name>OUT_6</name></connection>
<connection>
<GID>93</GID>
<name>IN_3</name></connection>
<connection>
<GID>61</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-26.5,130.5,-16.5</points>
<intersection>-26.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-26.5,144.5,-26.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<connection>
<GID>94</GID>
<name>IN_3</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-16.5,130.5,-16.5</points>
<connection>
<GID>113</GID>
<name>OUT_5</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-36,130,-17.5</points>
<intersection>-36 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-36,144.5,-36</points>
<connection>
<GID>63</GID>
<name>IN_3</name></connection>
<connection>
<GID>98</GID>
<name>IN_3</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-17.5,130,-17.5</points>
<connection>
<GID>113</GID>
<name>OUT_4</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-47,129.5,-18.5</points>
<intersection>-47 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-47,144.5,-47</points>
<connection>
<GID>64</GID>
<name>IN_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_3</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-18.5,129.5,-18.5</points>
<connection>
<GID>113</GID>
<name>OUT_3</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-58,129,-19.5</points>
<intersection>-58 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-58,144.5,-58</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-19.5,129,-19.5</points>
<connection>
<GID>113</GID>
<name>OUT_2</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-68.5,128.5,-20.5</points>
<intersection>-68.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-68.5,144.5,-68.5</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-20.5,128.5,-20.5</points>
<connection>
<GID>113</GID>
<name>OUT_1</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-79.5,128,-21.5</points>
<intersection>-79.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-21.5,128,-21.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-79.5,144.5,-79.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-27.5,127,-6.5</points>
<intersection>-27.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-6.5,144.5,-6.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-27.5,127,-27.5</points>
<connection>
<GID>114</GID>
<name>OUT_7</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-28.5,126.5,-17.5</points>
<intersection>-28.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-17.5,144.5,-17.5</points>
<connection>
<GID>61</GID>
<name>IN_2</name></connection>
<connection>
<GID>93</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-28.5,126.5,-28.5</points>
<connection>
<GID>114</GID>
<name>OUT_6</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-29.5,132,-29.5</points>
<connection>
<GID>114</GID>
<name>OUT_5</name></connection>
<intersection>132 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132,-29.5,132,-28.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-29.5 1</intersection>
<intersection>-28.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>132,-28.5,144.5,-28.5</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>132 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-38,126,-30.5</points>
<intersection>-38 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-38,144.5,-38</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-30.5,126,-30.5</points>
<connection>
<GID>114</GID>
<name>OUT_4</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-49,125.5,-31.5</points>
<intersection>-49 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-49,144.5,-49</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-31.5,125.5,-31.5</points>
<connection>
<GID>114</GID>
<name>OUT_3</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-60,125,-32.5</points>
<intersection>-60 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-60,144.5,-60</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-32.5,125,-32.5</points>
<connection>
<GID>114</GID>
<name>OUT_2</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-70.5,124.5,-33.5</points>
<intersection>-70.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-33.5,124.5,-33.5</points>
<connection>
<GID>114</GID>
<name>OUT_1</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-70.5,144.5,-70.5</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-81.5,127.5,-34.5</points>
<intersection>-81.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-81.5,144.5,-81.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-34.5,127.5,-34.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-41,123,-8.5</points>
<intersection>-41 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-8.5,144.5,-8.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-41,123,-41</points>
<connection>
<GID>58</GID>
<name>OUT_7</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-42,122.5,-19.5</points>
<intersection>-42 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-19.5,144.5,-19.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-42,122.5,-42</points>
<connection>
<GID>58</GID>
<name>OUT_6</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-43,122,-30.5</points>
<intersection>-43 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-30.5,144.5,-30.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-43,122,-43</points>
<connection>
<GID>58</GID>
<name>OUT_5</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-44,121.5,-40</points>
<intersection>-44 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-40,144.5,-40</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-44,121.5,-44</points>
<connection>
<GID>58</GID>
<name>OUT_4</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-51,121,-45</points>
<intersection>-51 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-51,144.5,-51</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-45,121,-45</points>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-62,120.5,-46</points>
<intersection>-62 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-62,144.5,-62</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-46,120.5,-46</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-72.5,120,-47</points>
<intersection>-72.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-72.5,144.5,-72.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-47,120,-47</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-83.5,119.5,-48</points>
<intersection>-83.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-48,119.5,-48</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-83.5,144.5,-83.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-54,118.5,-10.5</points>
<intersection>-54 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,-10.5,132,-10.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-54,118.5,-54</points>
<connection>
<GID>59</GID>
<name>OUT_7</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-55,118,-21.5</points>
<intersection>-55 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-21.5,144.5,-21.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-55,118,-55</points>
<connection>
<GID>59</GID>
<name>OUT_6</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-56,117.5,-32.5</points>
<intersection>-56 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-32.5,144.5,-32.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-56,117.5,-56</points>
<connection>
<GID>59</GID>
<name>OUT_5</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-42,144.5,-42</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>113.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113.5,-57,113.5,-42</points>
<connection>
<GID>59</GID>
<name>OUT_4</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-58,116.5,-53</points>
<intersection>-58 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-53,144.5,-53</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-58,116.5,-58</points>
<connection>
<GID>59</GID>
<name>OUT_3</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-64,116,-59</points>
<intersection>-64 1</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-64,144.5,-64</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-59,116,-59</points>
<connection>
<GID>59</GID>
<name>OUT_2</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-74.5,115.5,-60</points>
<intersection>-74.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-74.5,144.5,-74.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-60,115.5,-60</points>
<connection>
<GID>59</GID>
<name>OUT_1</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-36,156.5,-7.5</points>
<intersection>-36 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-7.5,156.5,-7.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-36,162,-36</points>
<connection>
<GID>70</GID>
<name>IN_7</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-37,156.5,-18.5</points>
<intersection>-37 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-18.5,156.5,-18.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-37,162,-37</points>
<connection>
<GID>70</GID>
<name>IN_6</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-38,156.5,-29.5</points>
<intersection>-38 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-29.5,156.5,-29.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-38,162,-38</points>
<connection>
<GID>70</GID>
<name>IN_5</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>138,-39,162,-39</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-50,156.5,-40</points>
<intersection>-50 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-50,156.5,-50</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-40,162,-40</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-61,156.5,-41</points>
<intersection>-61 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-61,156.5,-61</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-41,162,-41</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-71.5,156.5,-42</points>
<intersection>-71.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-71.5,156.5,-71.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156.5,-42,162,-42</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-82.5,156.5,-43</points>
<intersection>-82.5 2</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-43,162,-43</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-82.5,156.5,-82.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-85.5,115,-61</points>
<intersection>-85.5 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-85.5,144.5,-85.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-61,115,-61</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-66.5,105,-23.5</points>
<intersection>-66.5 10</intersection>
<intersection>-63 8</intersection>
<intersection>-50 7</intersection>
<intersection>-36.5 6</intersection>
<intersection>-23.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>105,-23.5,108.5,-23.5</points>
<connection>
<GID>113</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105,-36.5,108.5,-36.5</points>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>105,-50,108.5,-50</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>105,-63,108.5,-63</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>102,-66.5,105,-66.5</points>
<connection>
<GID>72</GID>
<name>CLK</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-77.5,136,0.5</points>
<connection>
<GID>69</GID>
<name>SEL_0</name></connection>
<connection>
<GID>66</GID>
<name>SEL_0</name></connection>
<connection>
<GID>65</GID>
<name>SEL_0</name></connection>
<connection>
<GID>64</GID>
<name>SEL_0</name></connection>
<connection>
<GID>63</GID>
<name>SEL_0</name></connection>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<connection>
<GID>61</GID>
<name>SEL_0</name></connection>
<connection>
<GID>60</GID>
<name>SEL_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,0.5,136,0.5</points>
<intersection>82.5 2</intersection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>82.5,-25.5,82.5,0.5</points>
<intersection>-25.5 3</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-25.5,82.5,-25.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>82.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-77.5,135,0</points>
<connection>
<GID>69</GID>
<name>SEL_1</name></connection>
<connection>
<GID>66</GID>
<name>SEL_1</name></connection>
<connection>
<GID>65</GID>
<name>SEL_1</name></connection>
<connection>
<GID>64</GID>
<name>SEL_1</name></connection>
<connection>
<GID>63</GID>
<name>SEL_1</name></connection>
<connection>
<GID>62</GID>
<name>SEL_1</name></connection>
<connection>
<GID>61</GID>
<name>SEL_1</name></connection>
<connection>
<GID>60</GID>
<name>SEL_1</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,0,135,0</points>
<intersection>82 2</intersection>
<intersection>135 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>82,-23.5,82,0</points>
<intersection>-23.5 3</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-23.5,82,-23.5</points>
<connection>
<GID>71</GID>
<name>OUT_1</name></connection>
<intersection>82 2</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-47,151,-7.5</points>
<intersection>-47 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-7.5,151,-7.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-47,162,-47</points>
<connection>
<GID>103</GID>
<name>IN_7</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-48,151,-18.5</points>
<intersection>-48 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-18.5,151,-18.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-48,162,-48</points>
<connection>
<GID>103</GID>
<name>IN_6</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-49,151,-29.5</points>
<intersection>-49 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-29.5,151,-29.5</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-49,162,-49</points>
<connection>
<GID>103</GID>
<name>IN_5</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-50,151,-39</points>
<intersection>-50 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-39,151,-39</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-50,162,-50</points>
<connection>
<GID>103</GID>
<name>IN_4</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-51,162,-51</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>151 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>151,-51,151,-50</points>
<intersection>-51 1</intersection>
<intersection>-50 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>150.5,-50,151,-50</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>151 2</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-61,151,-52</points>
<intersection>-61 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-61,151,-61</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-52,162,-52</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-71.5,151,-53</points>
<intersection>-71.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-71.5,151,-71.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-53,162,-53</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-82.5,151,-54</points>
<intersection>-82.5 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-54,162,-54</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>150.5,-82.5,151,-82.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-77.5,148.5,-1</points>
<connection>
<GID>102</GID>
<name>SEL_0</name></connection>
<connection>
<GID>101</GID>
<name>SEL_0</name></connection>
<connection>
<GID>100</GID>
<name>SEL_0</name></connection>
<connection>
<GID>99</GID>
<name>SEL_0</name></connection>
<connection>
<GID>98</GID>
<name>SEL_0</name></connection>
<connection>
<GID>94</GID>
<name>SEL_0</name></connection>
<connection>
<GID>93</GID>
<name>SEL_0</name></connection>
<connection>
<GID>87</GID>
<name>SEL_0</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-1,148.5,-1</points>
<intersection>83.5 2</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,-39.5,83.5,-1</points>
<intersection>-39.5 3</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-39.5,83.5,-39.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>83.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-77.5,147.5,-0.5</points>
<connection>
<GID>102</GID>
<name>SEL_1</name></connection>
<connection>
<GID>101</GID>
<name>SEL_1</name></connection>
<connection>
<GID>100</GID>
<name>SEL_1</name></connection>
<connection>
<GID>99</GID>
<name>SEL_1</name></connection>
<connection>
<GID>98</GID>
<name>SEL_1</name></connection>
<connection>
<GID>94</GID>
<name>SEL_1</name></connection>
<connection>
<GID>93</GID>
<name>SEL_1</name></connection>
<connection>
<GID>87</GID>
<name>SEL_1</name></connection>
<intersection>-0.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>83,-0.5,147.5,-0.5</points>
<intersection>83 16</intersection>
<intersection>147.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>83,-37.5,83,-0.5</points>
<intersection>-37.5 18</intersection>
<intersection>-0.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>81.5,-37.5,83,-37.5</points>
<connection>
<GID>78</GID>
<name>OUT_1</name></connection>
<intersection>83 16</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-54,104,-14.5</points>
<intersection>-54 6</intersection>
<intersection>-41 3</intersection>
<intersection>-33 4</intersection>
<intersection>-27.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-14.5,105.5,-14.5</points>
<connection>
<GID>113</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-27.5,105.5,-27.5</points>
<connection>
<GID>114</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-41,105.5,-41</points>
<connection>
<GID>58</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>97.5,-33,104,-33</points>
<connection>
<GID>105</GID>
<name>OUT_3</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104,-54,105.5,-54</points>
<connection>
<GID>59</GID>
<name>IN_7</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-55,103.5,-15.5</points>
<intersection>-55 6</intersection>
<intersection>-42 5</intersection>
<intersection>-35 2</intersection>
<intersection>-28.5 3</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-35,103.5,-35</points>
<connection>
<GID>105</GID>
<name>OUT_2</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,-28.5,105.5,-28.5</points>
<connection>
<GID>114</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103.5,-15.5,105.5,-15.5</points>
<connection>
<GID>113</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103.5,-42,105.5,-42</points>
<connection>
<GID>58</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103.5,-55,105.5,-55</points>
<connection>
<GID>59</GID>
<name>IN_6</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-56,103,-16.5</points>
<intersection>-56 6</intersection>
<intersection>-43 3</intersection>
<intersection>-37 2</intersection>
<intersection>-29.5 4</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-37,103,-37</points>
<connection>
<GID>105</GID>
<name>OUT_1</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,-43,105.5,-43</points>
<connection>
<GID>58</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103,-29.5,105.5,-29.5</points>
<connection>
<GID>114</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,-16.5,105.5,-16.5</points>
<connection>
<GID>113</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103,-56,105.5,-56</points>
<connection>
<GID>59</GID>
<name>IN_5</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-57,102.5,-17.5</points>
<intersection>-57 6</intersection>
<intersection>-44 3</intersection>
<intersection>-39 2</intersection>
<intersection>-30.5 4</intersection>
<intersection>-17.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-39,102.5,-39</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,-44,105.5,-44</points>
<connection>
<GID>58</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102.5,-30.5,105.5,-30.5</points>
<connection>
<GID>114</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102.5,-17.5,105.5,-17.5</points>
<connection>
<GID>113</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102.5,-57,105.5,-57</points>
<connection>
<GID>59</GID>
<name>IN_4</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-58,102,-18.5</points>
<intersection>-58 5</intersection>
<intersection>-45 2</intersection>
<intersection>-31.5 3</intersection>
<intersection>-18.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-45,105.5,-45</points>
<connection>
<GID>58</GID>
<name>IN_3</name></connection>
<connection>
<GID>106</GID>
<name>OUT_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,-31.5,105.5,-31.5</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102,-18.5,105.5,-18.5</points>
<connection>
<GID>113</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102,-58,105.5,-58</points>
<connection>
<GID>59</GID>
<name>IN_3</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-59,101.5,-19.5</points>
<intersection>-59 5</intersection>
<intersection>-47 2</intersection>
<intersection>-46 4</intersection>
<intersection>-32.5 3</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-19.5,105.5,-19.5</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-47,101.5,-47</points>
<connection>
<GID>106</GID>
<name>OUT_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-32.5,105.5,-32.5</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101.5,-46,105.5,-46</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101.5,-59,105.5,-59</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-60,101,-20.5</points>
<intersection>-60 5</intersection>
<intersection>-49 2</intersection>
<intersection>-47 4</intersection>
<intersection>-33.5 3</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-20.5,105.5,-20.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-49,101,-49</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-33.5,105.5,-33.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101,-47,105.5,-47</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101,-60,105.5,-60</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-61,100.5,-21.5</points>
<intersection>-61 5</intersection>
<intersection>-51 2</intersection>
<intersection>-48 4</intersection>
<intersection>-34.5 3</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-21.5,105.5,-21.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-51,100.5,-51</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>100.5,-34.5,105.5,-34.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>100.5,-48,105.5,-48</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>100.5,-61,105.5,-61</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-12.5,107.5,-4.5</points>
<intersection>-12.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-4.5,107.5,-4.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-12.5,108.5,-12.5</points>
<connection>
<GID>113</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-25.5,107.5,-3.5</points>
<intersection>-25.5 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-3.5,107.5,-3.5</points>
<connection>
<GID>108</GID>
<name>OUT_1</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-25.5,108.5,-25.5</points>
<connection>
<GID>114</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-39,107.5,-2.5</points>
<intersection>-39 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-2.5,107.5,-2.5</points>
<connection>
<GID>108</GID>
<name>OUT_2</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-39,108.5,-39</points>
<connection>
<GID>58</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-52,107.5,-1.5</points>
<intersection>-52 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-1.5,107.5,-1.5</points>
<connection>
<GID>108</GID>
<name>OUT_3</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-52,108.5,-52</points>
<connection>
<GID>59</GID>
<name>load</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-2.5,91.5,-2.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>91.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91.5,-2.5,91.5,-1.5</points>
<connection>
<GID>108</GID>
<name>ENABLE</name></connection>
<intersection>-2.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-18.5,96,-7.5</points>
<intersection>-18.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91,-7.5,96,-7.5</points>
<intersection>91 3</intersection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-18.5,96,-18.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91,-7.5,91,-4.5</points>
<intersection>-7.5 1</intersection>
<intersection>-4.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>91,-4.5,91.5,-4.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>91 3</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-16.5,96.5,-7</points>
<intersection>-16.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-7,96.5,-7</points>
<intersection>91.5 3</intersection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-16.5,96.5,-16.5</points>
<connection>
<GID>111</GID>
<name>OUT_1</name></connection>
<intersection>96.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-7,91.5,-3.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>10.5819,-1.68137,253.293,-129.863</PageViewport>
<gate>
<ID>196</ID>
<type>AA_INVERTER</type>
<position>70,-67.5</position>
<input>
<ID>IN_0</ID>268 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>94.5,-43</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>72,-75</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>72,-76.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AE_REGISTER8</type>
<position>99,-59</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>174 </input>
<input>
<ID>IN_2</ID>175 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_4</ID>177 </input>
<input>
<ID>IN_5</ID>178 </input>
<input>
<ID>IN_6</ID>179 </input>
<input>
<ID>IN_7</ID>180 </input>
<output>
<ID>OUT_0</ID>188 </output>
<output>
<ID>OUT_1</ID>187 </output>
<output>
<ID>OUT_2</ID>186 </output>
<output>
<ID>OUT_3</ID>185 </output>
<output>
<ID>OUT_4</ID>184 </output>
<output>
<ID>OUT_5</ID>183 </output>
<output>
<ID>OUT_6</ID>182 </output>
<output>
<ID>OUT_7</ID>181 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>267 </input>
<input>
<ID>count_enable</ID>203 </input>
<input>
<ID>count_up</ID>203 </input>
<input>
<ID>load</ID>269 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_REGISTER8</type>
<position>116,-59</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<input>
<ID>IN_2</ID>186 </input>
<input>
<ID>IN_3</ID>185 </input>
<input>
<ID>IN_4</ID>184 </input>
<input>
<ID>IN_5</ID>183 </input>
<input>
<ID>IN_6</ID>182 </input>
<input>
<ID>IN_7</ID>181 </input>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>217 </output>
<output>
<ID>OUT_2</ID>194 </output>
<output>
<ID>OUT_3</ID>193 </output>
<output>
<ID>OUT_4</ID>192 </output>
<output>
<ID>OUT_5</ID>191 </output>
<output>
<ID>OUT_6</ID>190 </output>
<output>
<ID>OUT_7</ID>189 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>202 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_REGISTER8</type>
<position>153,-76.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>256 </input>
<input>
<ID>IN_2</ID>257 </input>
<input>
<ID>IN_3</ID>258 </input>
<input>
<ID>IN_4</ID>259 </input>
<input>
<ID>IN_5</ID>254 </input>
<input>
<ID>IN_6</ID>261 </input>
<input>
<ID>IN_7</ID>260 </input>
<output>
<ID>OUT_0</ID>226 </output>
<output>
<ID>OUT_1</ID>225 </output>
<output>
<ID>OUT_2</ID>224 </output>
<output>
<ID>OUT_3</ID>223 </output>
<output>
<ID>OUT_4</ID>222 </output>
<output>
<ID>OUT_5</ID>221 </output>
<output>
<ID>OUT_6</ID>220 </output>
<output>
<ID>OUT_7</ID>219 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>216 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_RAM_8x8</type>
<position>131,-58.5</position>
<input>
<ID>ADDRESS_0</ID>218 </input>
<input>
<ID>ADDRESS_1</ID>217 </input>
<input>
<ID>ADDRESS_2</ID>194 </input>
<input>
<ID>ADDRESS_3</ID>193 </input>
<input>
<ID>ADDRESS_4</ID>192 </input>
<input>
<ID>ADDRESS_5</ID>191 </input>
<input>
<ID>ADDRESS_6</ID>190 </input>
<input>
<ID>ADDRESS_7</ID>189 </input>
<input>
<ID>DATA_IN_0</ID>262 </input>
<input>
<ID>DATA_IN_1</ID>242 </input>
<input>
<ID>DATA_IN_2</ID>245 </input>
<input>
<ID>DATA_IN_3</ID>246 </input>
<input>
<ID>DATA_IN_4</ID>247 </input>
<input>
<ID>DATA_IN_5</ID>251 </input>
<input>
<ID>DATA_IN_6</ID>252 </input>
<input>
<ID>DATA_IN_7</ID>253 </input>
<output>
<ID>DATA_OUT_0</ID>262 </output>
<output>
<ID>DATA_OUT_1</ID>242 </output>
<output>
<ID>DATA_OUT_2</ID>245 </output>
<output>
<ID>DATA_OUT_3</ID>246 </output>
<output>
<ID>DATA_OUT_4</ID>247 </output>
<output>
<ID>DATA_OUT_5</ID>251 </output>
<output>
<ID>DATA_OUT_6</ID>252 </output>
<output>
<ID>DATA_OUT_7</ID>253 </output>
<input>
<ID>ENABLE_0</ID>241 </input>
<input>
<ID>write_enable</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 170</lparam>
<lparam>Address:1 187</lparam>
<lparam>Address:2 204</lparam>
<lparam>Address:3 221</lparam></gate>
<gate>
<ID>127</ID>
<type>AE_REGISTER8</type>
<position>169,-76.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>225 </input>
<input>
<ID>IN_2</ID>224 </input>
<input>
<ID>IN_3</ID>223 </input>
<input>
<ID>IN_4</ID>222 </input>
<input>
<ID>IN_5</ID>221 </input>
<input>
<ID>IN_6</ID>220 </input>
<input>
<ID>IN_7</ID>219 </input>
<output>
<ID>OUT_0</ID>236 </output>
<output>
<ID>OUT_1</ID>237 </output>
<input>
<ID>clear</ID>239 </input>
<input>
<ID>clock</ID>238 </input>
<input>
<ID>load</ID>227 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>131</ID>
<type>DD_KEYPAD_HEX</type>
<position>79.5,-65</position>
<output>
<ID>OUT_0</ID>173 </output>
<output>
<ID>OUT_1</ID>174 </output>
<output>
<ID>OUT_2</ID>175 </output>
<output>
<ID>OUT_3</ID>176 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>133</ID>
<type>DD_KEYPAD_HEX</type>
<position>79.5,-53</position>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>178 </output>
<output>
<ID>OUT_2</ID>179 </output>
<output>
<ID>OUT_3</ID>180 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>135</ID>
<type>BB_CLOCK</type>
<position>68,-90.5</position>
<output>
<ID>CLK</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>97,-40</position>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>84.5,-42</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>84.5,-39.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>110,-42.5</position>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>98,-87.5</position>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>92.5,-84.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>149,-69</position>
<output>
<ID>OUT_0</ID>216 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>94,-51</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>110.5,-51</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>131,-50</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>153,-66</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>166,-68.5</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>169</ID>
<type>BE_ROM_8x8</type>
<position>184,-76</position>
<input>
<ID>ADDRESS_0</ID>236 </input>
<input>
<ID>ADDRESS_1</ID>237 </input>
<input>
<ID>ENABLE_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>141,-56</position>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>141,-59</position>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>147.5,-55.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>148,-58.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>145,-76</position>
<input>
<ID>ENABLE_0</ID>241 </input>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>245 </input>
<input>
<ID>IN_3</ID>246 </input>
<input>
<ID>IN_4</ID>247 </input>
<input>
<ID>IN_5</ID>251 </input>
<input>
<ID>IN_6</ID>252 </input>
<input>
<ID>IN_7</ID>253 </input>
<output>
<ID>OUT_0</ID>255 </output>
<output>
<ID>OUT_1</ID>256 </output>
<output>
<ID>OUT_2</ID>257 </output>
<output>
<ID>OUT_3</ID>258 </output>
<output>
<ID>OUT_4</ID>259 </output>
<output>
<ID>OUT_5</ID>254 </output>
<output>
<ID>OUT_6</ID>261 </output>
<output>
<ID>OUT_7</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>178</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>124,-76</position>
<input>
<ID>ENABLE_0</ID>240 </input>
<output>
<ID>OUT_0</ID>262 </output>
<output>
<ID>OUT_1</ID>242 </output>
<output>
<ID>OUT_2</ID>245 </output>
<output>
<ID>OUT_3</ID>246 </output>
<output>
<ID>OUT_4</ID>247 </output>
<output>
<ID>OUT_5</ID>251 </output>
<output>
<ID>OUT_6</ID>252 </output>
<output>
<ID>OUT_7</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>170.5,-68</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>193,-76.5</position>
<output>
<ID>OUT_0</ID>264 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>194.5,-73.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_AND2</type>
<position>94,-72</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>79.5,-89.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>74,-86.5</position>
<output>
<ID>OUT_0</ID>266 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>65,-73</position>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-59,126,-59</points>
<connection>
<GID>119</GID>
<name>OUT_3</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-60,126,-60</points>
<connection>
<GID>119</GID>
<name>OUT_2</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-53,115,-42.5</points>
<connection>
<GID>119</GID>
<name>load</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-42.5,115,-42.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-53,99,-40</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>count_enable</name></connection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99,-52,100,-52</points>
<intersection>99 0</intersection>
<intersection>100 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100,-53,100,-52</points>
<connection>
<GID>117</GID>
<name>count_up</name></connection>
<intersection>-52 2</intersection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>151,-69,152,-69</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>152 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>152,-70.5,152,-69</points>
<connection>
<GID>123</GID>
<name>load</name></connection>
<intersection>-69 2</intersection></vsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-61,126,-61</points>
<connection>
<GID>119</GID>
<name>OUT_1</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-62,126,-62</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-72.5,165,-72.5</points>
<connection>
<GID>123</GID>
<name>OUT_7</name></connection>
<connection>
<GID>127</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-73.5,165,-73.5</points>
<connection>
<GID>123</GID>
<name>OUT_6</name></connection>
<connection>
<GID>127</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-74.5,165,-74.5</points>
<connection>
<GID>123</GID>
<name>OUT_5</name></connection>
<connection>
<GID>127</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-75.5,165,-75.5</points>
<connection>
<GID>123</GID>
<name>OUT_4</name></connection>
<connection>
<GID>127</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-76.5,165,-76.5</points>
<connection>
<GID>123</GID>
<name>OUT_3</name></connection>
<connection>
<GID>127</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-77.5,165,-77.5</points>
<connection>
<GID>123</GID>
<name>OUT_2</name></connection>
<connection>
<GID>127</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-78.5,165,-78.5</points>
<connection>
<GID>123</GID>
<name>OUT_1</name></connection>
<connection>
<GID>127</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-79.5,165,-79.5</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-70.5,168,-68.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<connection>
<GID>127</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173,-79.5,179,-79.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<connection>
<GID>169</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>173,-78.5,179,-78.5</points>
<connection>
<GID>127</GID>
<name>OUT_1</name></connection>
<connection>
<GID>169</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-89.5,115,-64</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-89.5,168,-89.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>85 6</intersection>
<intersection>115 0</intersection>
<intersection>152 5</intersection>
<intersection>168 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>168,-89.5,168,-81.5</points>
<connection>
<GID>127</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>152,-89.5,152,-81.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>85,-89.5,85,-71</points>
<intersection>-89.5 1</intersection>
<intersection>-71 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>85,-71,91,-71</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>85 6</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-87.5,100,-64</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,-87.5,170,-87.5</points>
<intersection>100 0</intersection>
<intersection>117 3</intersection>
<intersection>154 7</intersection>
<intersection>170 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>117,-87.5,117,-64</points>
<connection>
<GID>119</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>170,-87.5,170,-81.5</points>
<connection>
<GID>127</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>154,-87.5,154,-81.5</points>
<connection>
<GID>123</GID>
<name>clear</name></connection>
<intersection>-87.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-56,139,-56</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>136 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>136,-71,136,-56</points>
<connection>
<GID>125</GID>
<name>write_enable</name></connection>
<intersection>-71 4</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,-71,136,-71</points>
<connection>
<GID>178</GID>
<name>ENABLE_0</name></connection>
<intersection>136 3</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,-59,139,-59</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>ENABLE_0</name></connection>
<intersection>139 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>139,-71,139,-59</points>
<intersection>-71 6</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>139,-71,145,-71</points>
<connection>
<GID>177</GID>
<name>ENABLE_0</name></connection>
<intersection>139 5</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-78.5,143,-78.5</points>
<connection>
<GID>178</GID>
<name>OUT_1</name></connection>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>133.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>133.5,-78.5,133.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-77.5,143,-77.5</points>
<connection>
<GID>178</GID>
<name>OUT_2</name></connection>
<connection>
<GID>177</GID>
<name>IN_2</name></connection>
<intersection>132.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132.5,-77.5,132.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_2</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-76.5,143,-76.5</points>
<connection>
<GID>178</GID>
<name>OUT_3</name></connection>
<connection>
<GID>177</GID>
<name>IN_3</name></connection>
<intersection>131.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>131.5,-76.5,131.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_3</name></connection>
<intersection>-76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-75.5,143,-75.5</points>
<connection>
<GID>178</GID>
<name>OUT_4</name></connection>
<connection>
<GID>177</GID>
<name>IN_4</name></connection>
<intersection>130.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130.5,-75.5,130.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_4</name></connection>
<intersection>-75.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-74.5,143,-74.5</points>
<connection>
<GID>178</GID>
<name>OUT_5</name></connection>
<connection>
<GID>177</GID>
<name>IN_5</name></connection>
<intersection>129.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>129.5,-74.5,129.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_5</name></connection>
<intersection>-74.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-73.5,143,-73.5</points>
<connection>
<GID>178</GID>
<name>OUT_6</name></connection>
<connection>
<GID>177</GID>
<name>IN_6</name></connection>
<intersection>128.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-73.5,128.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_6</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-72.5,143,-72.5</points>
<connection>
<GID>178</GID>
<name>OUT_7</name></connection>
<connection>
<GID>177</GID>
<name>IN_7</name></connection>
<intersection>127.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127.5,-72.5,127.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_7</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-74.5,149,-74.5</points>
<connection>
<GID>123</GID>
<name>IN_5</name></connection>
<connection>
<GID>177</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-79.5,149,-79.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-78.5,149,-78.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<connection>
<GID>177</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-77.5,149,-77.5</points>
<connection>
<GID>123</GID>
<name>IN_2</name></connection>
<connection>
<GID>177</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-76.5,149,-76.5</points>
<connection>
<GID>123</GID>
<name>IN_3</name></connection>
<connection>
<GID>177</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-75.5,149,-75.5</points>
<connection>
<GID>123</GID>
<name>IN_4</name></connection>
<connection>
<GID>177</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-72.5,149,-72.5</points>
<connection>
<GID>123</GID>
<name>IN_7</name></connection>
<connection>
<GID>177</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-73.5,149,-73.5</points>
<connection>
<GID>123</GID>
<name>IN_6</name></connection>
<connection>
<GID>177</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-79.5,143,-79.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>134.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-79.5,134.5,-65.5</points>
<connection>
<GID>125</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>DATA_IN_0</name></connection>
<intersection>-79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189,-76.5,191,-76.5</points>
<connection>
<GID>169</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-90.5,76.5,-90.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-88.5,76.5,-86.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-86.5,76.5,-86.5</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-72,98,-64</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-72,98,-72</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-73,91,-73</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>70 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>70,-73,70,-70.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-73 1</intersection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-53,98,-45</points>
<connection>
<GID>117</GID>
<name>load</name></connection>
<intersection>-45 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-64.5,70,-45</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-45,98,-45</points>
<intersection>70 1</intersection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-68,89.5,-62</points>
<intersection>-68 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-62,95,-62</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-68,89.5,-68</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-66,89.5,-61</points>
<intersection>-66 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-61,95,-61</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-66,89.5,-66</points>
<connection>
<GID>131</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-64,89.5,-60</points>
<intersection>-64 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-60,95,-60</points>
<connection>
<GID>117</GID>
<name>IN_2</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-64,89.5,-64</points>
<connection>
<GID>131</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-62,89.5,-59</points>
<intersection>-62 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-59,95,-59</points>
<connection>
<GID>117</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-62,89.5,-62</points>
<connection>
<GID>131</GID>
<name>OUT_3</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-58,89.5,-56</points>
<intersection>-58 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-58,95,-58</points>
<connection>
<GID>117</GID>
<name>IN_4</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-56,89.5,-56</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-57,89.5,-54</points>
<intersection>-57 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-57,95,-57</points>
<connection>
<GID>117</GID>
<name>IN_5</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-54,89.5,-54</points>
<connection>
<GID>133</GID>
<name>OUT_1</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-56,89.5,-52</points>
<intersection>-56 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-56,95,-56</points>
<connection>
<GID>117</GID>
<name>IN_6</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-52,89.5,-52</points>
<connection>
<GID>133</GID>
<name>OUT_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-55,95,-55</points>
<connection>
<GID>117</GID>
<name>IN_7</name></connection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-55,84.5,-50</points>
<connection>
<GID>133</GID>
<name>OUT_3</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-55,112,-55</points>
<connection>
<GID>119</GID>
<name>IN_7</name></connection>
<connection>
<GID>117</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-56,112,-56</points>
<connection>
<GID>119</GID>
<name>IN_6</name></connection>
<connection>
<GID>117</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-57,112,-57</points>
<connection>
<GID>119</GID>
<name>IN_5</name></connection>
<connection>
<GID>117</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-58,112,-58</points>
<connection>
<GID>119</GID>
<name>IN_4</name></connection>
<connection>
<GID>117</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-59,112,-59</points>
<connection>
<GID>119</GID>
<name>IN_3</name></connection>
<connection>
<GID>117</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-60,112,-60</points>
<connection>
<GID>119</GID>
<name>IN_2</name></connection>
<connection>
<GID>117</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-61,112,-61</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<connection>
<GID>117</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-62,112,-62</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-55,126,-55</points>
<connection>
<GID>119</GID>
<name>OUT_7</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-56,126,-56</points>
<connection>
<GID>119</GID>
<name>OUT_6</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-57,126,-57</points>
<connection>
<GID>119</GID>
<name>OUT_5</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-58,126,-58</points>
<connection>
<GID>119</GID>
<name>OUT_4</name></connection>
<connection>
<GID>125</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-153.642,84.6798,497.642,-259.278</PageViewport>
<gate>
<ID>1484</ID>
<type>AA_LABEL</type>
<position>125,-71</position>
<gparam>LABEL_TEXT Skip to page 5</gparam>
<gparam>TEXT_HEIGHT 20</gparam>
<gparam>angle 0.0</gparam></gate></page 3>
<page 4>
<PageViewport>-92.75,54.4618,284.75,-144.904</PageViewport>
<gate>
<ID>386</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-93</position>
<output>
<ID>OUT_0</ID>545 </output>
<output>
<ID>OUT_1</ID>547 </output>
<output>
<ID>OUT_2</ID>549 </output>
<output>
<ID>OUT_3</ID>551 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>387</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-117</position>
<output>
<ID>OUT_0</ID>544 </output>
<output>
<ID>OUT_1</ID>546 </output>
<output>
<ID>OUT_2</ID>548 </output>
<output>
<ID>OUT_3</ID>550 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>-35.5,-106</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>389</ID>
<type>AA_LABEL</type>
<position>-36,-80</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>AA_LABEL</type>
<position>-36,-92.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>AA_LABEL</type>
<position>-36,-117.5</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>BA_DECODER_2x4</type>
<position>5.5,-71</position>
<input>
<ID>ENABLE</ID>560 </input>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>562 </output>
<output>
<ID>OUT_1</ID>563 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_TOGGLE</type>
<position>0.5,-69.5</position>
<output>
<ID>OUT_0</ID>560 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_TOGGLE</type>
<position>-4,-72.5</position>
<output>
<ID>OUT_0</ID>561 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_LABEL</type>
<position>1,-66.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_LABEL</type>
<position>-10.5,-72</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,-106.5</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>574 </input>
<input>
<ID>IN_2</ID>575 </input>
<input>
<ID>IN_3</ID>576 </input>
<input>
<ID>IN_B_0</ID>565 </input>
<input>
<ID>IN_B_1</ID>566 </input>
<input>
<ID>IN_B_2</ID>567 </input>
<input>
<ID>IN_B_3</ID>568 </input>
<output>
<ID>OUT_0</ID>597 </output>
<output>
<ID>OUT_1</ID>598 </output>
<output>
<ID>OUT_2</ID>599 </output>
<output>
<ID>OUT_3</ID>600 </output>
<output>
<ID>carry_out</ID>564 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>398</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31.5,-122.5</position>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>578 </input>
<input>
<ID>IN_2</ID>579 </input>
<input>
<ID>IN_3</ID>580 </input>
<input>
<ID>IN_B_0</ID>569 </input>
<input>
<ID>IN_B_1</ID>570 </input>
<input>
<ID>IN_B_2</ID>571 </input>
<input>
<ID>IN_B_3</ID>572 </input>
<output>
<ID>OUT_0</ID>601 </output>
<output>
<ID>OUT_1</ID>602 </output>
<output>
<ID>OUT_2</ID>603 </output>
<output>
<ID>OUT_3</ID>604 </output>
<input>
<ID>carry_in</ID>564 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>399</ID>
<type>AA_LABEL</type>
<position>39,-99</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>39.5,-127.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_LABEL</type>
<position>25,-100</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>AA_LABEL</type>
<position>25.5,-106.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AA_LABEL</type>
<position>25,-116</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>AA_LABEL</type>
<position>26,-123</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>27,-96</position>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>32,-92.5</position>
<input>
<ID>IN_0</ID>584 </input>
<input>
<ID>IN_1</ID>583 </input>
<output>
<ID>OUT</ID>606 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>27,-89</position>
<input>
<ID>IN_0</ID>586 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>32,-85.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>587 </input>
<output>
<ID>OUT</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>27,-82</position>
<input>
<ID>IN_0</ID>590 </input>
<input>
<ID>IN_1</ID>589 </input>
<output>
<ID>OUT</ID>609 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>32,-78.5</position>
<input>
<ID>IN_0</ID>592 </input>
<input>
<ID>IN_1</ID>591 </input>
<output>
<ID>OUT</ID>610 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_AND2</type>
<position>27,-75</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>593 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_AND2</type>
<position>32,-71.5</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>595 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>413</ID>
<type>AA_MUX_2x1</type>
<position>57,-83</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>612 </input>
<output>
<ID>OUT</ID>620 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>AA_MUX_2x1</type>
<position>57,-88</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>611 </input>
<output>
<ID>OUT</ID>619 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_MUX_2x1</type>
<position>57,-93</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>610 </input>
<output>
<ID>OUT</ID>618 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_MUX_2x1</type>
<position>57,-98</position>
<input>
<ID>IN_0</ID>601 </input>
<input>
<ID>IN_1</ID>609 </input>
<output>
<ID>OUT</ID>617 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>AA_MUX_2x1</type>
<position>57,-103</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>608 </input>
<output>
<ID>OUT</ID>616 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_MUX_2x1</type>
<position>57,-108</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>615 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_MUX_2x1</type>
<position>57,-113</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>614 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_MUX_2x1</type>
<position>57,-118</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>605 </input>
<output>
<ID>OUT</ID>613 </output>
<input>
<ID>SEL_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>79.5,-100</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>614 </input>
<input>
<ID>IN_2</ID>615 </input>
<input>
<ID>IN_3</ID>616 </input>
<input>
<ID>IN_4</ID>617 </input>
<input>
<ID>IN_5</ID>618 </input>
<input>
<ID>IN_6</ID>619 </input>
<input>
<ID>IN_7</ID>620 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 54</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>422</ID>
<type>AA_LABEL</type>
<position>57,-121.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>58,-79</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>424</ID>
<type>GA_LED</type>
<position>71,-110</position>
<input>
<ID>N_in2</ID>620 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>425</ID>
<type>GA_LED</type>
<position>73.5,-110</position>
<input>
<ID>N_in2</ID>619 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>426</ID>
<type>GA_LED</type>
<position>76,-110</position>
<input>
<ID>N_in2</ID>618 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>427</ID>
<type>GA_LED</type>
<position>78.5,-110</position>
<input>
<ID>N_in2</ID>617 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>428</ID>
<type>GA_LED</type>
<position>81,-110</position>
<input>
<ID>N_in2</ID>616 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>429</ID>
<type>GA_LED</type>
<position>83.5,-110</position>
<input>
<ID>N_in2</ID>615 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>430</ID>
<type>GA_LED</type>
<position>86,-110</position>
<input>
<ID>N_in2</ID>614 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>431</ID>
<type>GA_LED</type>
<position>88.5,-110</position>
<input>
<ID>N_in2</ID>613 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>88.5,-112</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AA_LABEL</type>
<position>86,-112</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>83.5,-112</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>81,-112</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>78.5,-112</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AA_LABEL</type>
<position>76,-112</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>73.5,-112</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>71,-112</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>207,-63.5</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>AA_LABEL</type>
<position>207,-74.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>AE_REGISTER8</type>
<position>150,-74.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>644 </output>
<output>
<ID>OUT_1</ID>643 </output>
<output>
<ID>OUT_2</ID>642 </output>
<output>
<ID>OUT_3</ID>641 </output>
<output>
<ID>OUT_4</ID>640 </output>
<output>
<ID>OUT_5</ID>639 </output>
<output>
<ID>OUT_6</ID>638 </output>
<output>
<ID>OUT_7</ID>637 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>684 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>443</ID>
<type>AE_REGISTER8</type>
<position>150,-87.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>660 </output>
<output>
<ID>OUT_1</ID>651 </output>
<output>
<ID>OUT_2</ID>650 </output>
<output>
<ID>OUT_3</ID>649 </output>
<output>
<ID>OUT_4</ID>648 </output>
<output>
<ID>OUT_5</ID>647 </output>
<output>
<ID>OUT_6</ID>646 </output>
<output>
<ID>OUT_7</ID>645 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>685 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>444</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-37</position>
<input>
<ID>IN_0</ID>645 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>621 </input>
<output>
<ID>OUT</ID>652 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>445</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-48</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>638 </input>
<input>
<ID>IN_2</ID>630 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>653 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>446</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-59</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>639 </input>
<input>
<ID>IN_2</ID>631 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT</ID>654 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>447</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-68.5</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>640 </input>
<input>
<ID>IN_2</ID>632 </input>
<input>
<ID>IN_3</ID>624 </input>
<output>
<ID>OUT</ID>655 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-79.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>641 </input>
<input>
<ID>IN_2</ID>633 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT</ID>656 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-90.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>642 </input>
<input>
<ID>IN_2</ID>634 </input>
<input>
<ID>IN_3</ID>626 </input>
<output>
<ID>OUT</ID>657 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>450</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-101</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>643 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>658 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>451</ID>
<type>AE_MUX_4x1</type>
<position>175.5,-112</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>644 </input>
<input>
<ID>IN_2</ID>636 </input>
<input>
<ID>IN_3</ID>628 </input>
<output>
<ID>OUT</ID>659 </output>
<input>
<ID>SEL_0</ID>662 </input>
<input>
<ID>SEL_1</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>452</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>207.5,-69.5</position>
<input>
<ID>IN_0</ID>659 </input>
<input>
<ID>IN_1</ID>658 </input>
<input>
<ID>IN_2</ID>657 </input>
<input>
<ID>IN_3</ID>656 </input>
<input>
<ID>IN_4</ID>655 </input>
<input>
<ID>IN_5</ID>654 </input>
<input>
<ID>IN_6</ID>653 </input>
<input>
<ID>IN_7</ID>652 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>453</ID>
<type>DD_KEYPAD_HEX</type>
<position>117,-52</position>
<output>
<ID>OUT_0</ID>662 </output>
<output>
<ID>OUT_1</ID>663 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>454</ID>
<type>BB_CLOCK</type>
<position>138.5,-96</position>
<output>
<ID>CLK</ID>661 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>151,-41</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>151,-54</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_LABEL</type>
<position>151,-67.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AA_LABEL</type>
<position>151,-80.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>459</ID>
<type>AA_LABEL</type>
<position>115.5,-45</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>460</ID>
<type>DD_KEYPAD_HEX</type>
<position>117,-66</position>
<output>
<ID>OUT_0</ID>672 </output>
<output>
<ID>OUT_1</ID>673 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_MUX_4x1</type>
<position>188,-37</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>629 </input>
<input>
<ID>IN_3</ID>621 </input>
<output>
<ID>OUT</ID>664 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_MUX_4x1</type>
<position>188,-48</position>
<input>
<ID>IN_0</ID>646 </input>
<input>
<ID>IN_1</ID>638 </input>
<input>
<ID>IN_2</ID>630 </input>
<input>
<ID>IN_3</ID>622 </input>
<output>
<ID>OUT</ID>665 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_MUX_4x1</type>
<position>188,-59</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>639 </input>
<input>
<ID>IN_2</ID>631 </input>
<input>
<ID>IN_3</ID>623 </input>
<output>
<ID>OUT</ID>666 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_MUX_4x1</type>
<position>188,-68.5</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>640 </input>
<input>
<ID>IN_2</ID>632 </input>
<input>
<ID>IN_3</ID>624 </input>
<output>
<ID>OUT</ID>667 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>465</ID>
<type>AE_MUX_4x1</type>
<position>188,-79.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>641 </input>
<input>
<ID>IN_2</ID>633 </input>
<input>
<ID>IN_3</ID>625 </input>
<output>
<ID>OUT</ID>668 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>466</ID>
<type>AE_MUX_4x1</type>
<position>188,-90.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>642 </input>
<input>
<ID>IN_2</ID>634 </input>
<input>
<ID>IN_3</ID>626 </input>
<output>
<ID>OUT</ID>669 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_MUX_4x1</type>
<position>188,-101</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>643 </input>
<input>
<ID>IN_2</ID>635 </input>
<input>
<ID>IN_3</ID>627 </input>
<output>
<ID>OUT</ID>670 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>468</ID>
<type>AE_MUX_4x1</type>
<position>188,-112</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>644 </input>
<input>
<ID>IN_2</ID>636 </input>
<input>
<ID>IN_3</ID>628 </input>
<output>
<ID>OUT</ID>671 </output>
<input>
<ID>SEL_0</ID>672 </input>
<input>
<ID>SEL_1</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>469</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>207.5,-80.5</position>
<input>
<ID>IN_0</ID>671 </input>
<input>
<ID>IN_1</ID>670 </input>
<input>
<ID>IN_2</ID>669 </input>
<input>
<ID>IN_3</ID>668 </input>
<input>
<ID>IN_4</ID>667 </input>
<input>
<ID>IN_5</ID>666 </input>
<input>
<ID>IN_6</ID>665 </input>
<input>
<ID>IN_7</ID>664 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_LABEL</type>
<position>115.5,-59</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>DD_KEYPAD_HEX</type>
<position>133,-65.5</position>
<output>
<ID>OUT_0</ID>677 </output>
<output>
<ID>OUT_1</ID>676 </output>
<output>
<ID>OUT_2</ID>675 </output>
<output>
<ID>OUT_3</ID>674 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>472</ID>
<type>DD_KEYPAD_HEX</type>
<position>133,-77.5</position>
<output>
<ID>OUT_0</ID>681 </output>
<output>
<ID>OUT_1</ID>680 </output>
<output>
<ID>OUT_2</ID>679 </output>
<output>
<ID>OUT_3</ID>678 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>473</ID>
<type>AA_LABEL</type>
<position>133,-58.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>BA_DECODER_2x4</type>
<position>135,-32.5</position>
<input>
<ID>ENABLE</ID>686 </input>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>688 </input>
<output>
<ID>OUT_0</ID>682 </output>
<output>
<ID>OUT_1</ID>683 </output>
<output>
<ID>OUT_2</ID>684 </output>
<output>
<ID>OUT_3</ID>685 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_TOGGLE</type>
<position>129,-32</position>
<output>
<ID>OUT_0</ID>686 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>476</ID>
<type>AA_LABEL</type>
<position>126.5,-30.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>477</ID>
<type>DD_KEYPAD_HEX</type>
<position>130,-45</position>
<output>
<ID>OUT_0</ID>687 </output>
<output>
<ID>OUT_1</ID>688 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>130.5,-38</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>AE_REGISTER8</type>
<position>150,-48</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>628 </output>
<output>
<ID>OUT_1</ID>627 </output>
<output>
<ID>OUT_2</ID>626 </output>
<output>
<ID>OUT_3</ID>625 </output>
<output>
<ID>OUT_4</ID>624 </output>
<output>
<ID>OUT_5</ID>623 </output>
<output>
<ID>OUT_6</ID>622 </output>
<output>
<ID>OUT_7</ID>621 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>682 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>480</ID>
<type>AE_REGISTER8</type>
<position>150,-61</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<input>
<ID>IN_2</ID>679 </input>
<input>
<ID>IN_3</ID>678 </input>
<input>
<ID>IN_4</ID>677 </input>
<input>
<ID>IN_5</ID>676 </input>
<input>
<ID>IN_6</ID>675 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT_0</ID>636 </output>
<output>
<ID>OUT_1</ID>635 </output>
<output>
<ID>OUT_2</ID>634 </output>
<output>
<ID>OUT_3</ID>633 </output>
<output>
<ID>OUT_4</ID>632 </output>
<output>
<ID>OUT_5</ID>631 </output>
<output>
<ID>OUT_6</ID>630 </output>
<output>
<ID>OUT_7</ID>629 </output>
<input>
<ID>clock</ID>661 </input>
<input>
<ID>load</ID>683 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>481</ID>
<type>AA_LABEL</type>
<position>160.5,-23.5</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>483</ID>
<type>AA_LABEL</type>
<position>19.5,-37</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>485</ID>
<type>AA_LABEL</type>
<position>96,37.5</position>
<gparam>LABEL_TEXT Last update before starting to connect the pieces</gparam>
<gparam>TEXT_HEIGHT 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>87.5,20.5</position>
<gparam>LABEL_TEXT Check page 6</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>AA_INVERTER</type>
<position>-34,-23.5</position>
<input>
<ID>IN_0</ID>542 </input>
<output>
<ID>OUT_0</ID>543 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_TOGGLE</type>
<position>-9.5,1</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_LABEL</type>
<position>-32,-31</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>AA_LABEL</type>
<position>-32,-32.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AE_REGISTER8</type>
<position>-5,-15</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>481 </input>
<input>
<ID>IN_2</ID>482 </input>
<input>
<ID>IN_3</ID>483 </input>
<input>
<ID>IN_4</ID>484 </input>
<input>
<ID>IN_5</ID>485 </input>
<input>
<ID>IN_6</ID>486 </input>
<input>
<ID>IN_7</ID>487 </input>
<output>
<ID>OUT_0</ID>495 </output>
<output>
<ID>OUT_1</ID>494 </output>
<output>
<ID>OUT_2</ID>493 </output>
<output>
<ID>OUT_3</ID>492 </output>
<output>
<ID>OUT_4</ID>491 </output>
<output>
<ID>OUT_5</ID>490 </output>
<output>
<ID>OUT_6</ID>489 </output>
<output>
<ID>OUT_7</ID>488 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>541 </input>
<input>
<ID>count_enable</ID>503 </input>
<input>
<ID>count_up</ID>503 </input>
<input>
<ID>load</ID>543 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>348</ID>
<type>AE_REGISTER8</type>
<position>12,-15</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>494 </input>
<input>
<ID>IN_2</ID>493 </input>
<input>
<ID>IN_3</ID>492 </input>
<input>
<ID>IN_4</ID>491 </input>
<input>
<ID>IN_5</ID>490 </input>
<input>
<ID>IN_6</ID>489 </input>
<input>
<ID>IN_7</ID>488 </input>
<output>
<ID>OUT_0</ID>506 </output>
<output>
<ID>OUT_1</ID>505 </output>
<output>
<ID>OUT_2</ID>501 </output>
<output>
<ID>OUT_3</ID>500 </output>
<output>
<ID>OUT_4</ID>499 </output>
<output>
<ID>OUT_5</ID>498 </output>
<output>
<ID>OUT_6</ID>497 </output>
<output>
<ID>OUT_7</ID>496 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>502 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>349</ID>
<type>AE_REGISTER8</type>
<position>49,-32.5</position>
<input>
<ID>IN_0</ID>530 </input>
<input>
<ID>IN_1</ID>531 </input>
<input>
<ID>IN_2</ID>532 </input>
<input>
<ID>IN_3</ID>533 </input>
<input>
<ID>IN_4</ID>534 </input>
<input>
<ID>IN_5</ID>529 </input>
<input>
<ID>IN_6</ID>536 </input>
<input>
<ID>IN_7</ID>535 </input>
<output>
<ID>OUT_0</ID>514 </output>
<output>
<ID>OUT_1</ID>513 </output>
<output>
<ID>OUT_2</ID>512 </output>
<output>
<ID>OUT_3</ID>511 </output>
<output>
<ID>OUT_4</ID>510 </output>
<output>
<ID>OUT_5</ID>509 </output>
<output>
<ID>OUT_6</ID>508 </output>
<output>
<ID>OUT_7</ID>507 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>504 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_RAM_8x8</type>
<position>27,-14.5</position>
<input>
<ID>ADDRESS_0</ID>506 </input>
<input>
<ID>ADDRESS_1</ID>505 </input>
<input>
<ID>ADDRESS_2</ID>501 </input>
<input>
<ID>ADDRESS_3</ID>500 </input>
<input>
<ID>ADDRESS_4</ID>499 </input>
<input>
<ID>ADDRESS_5</ID>498 </input>
<input>
<ID>ADDRESS_6</ID>497 </input>
<input>
<ID>ADDRESS_7</ID>496 </input>
<input>
<ID>DATA_IN_0</ID>537 </input>
<input>
<ID>DATA_IN_1</ID>522 </input>
<input>
<ID>DATA_IN_2</ID>523 </input>
<input>
<ID>DATA_IN_3</ID>524 </input>
<input>
<ID>DATA_IN_4</ID>525 </input>
<input>
<ID>DATA_IN_5</ID>526 </input>
<input>
<ID>DATA_IN_6</ID>527 </input>
<input>
<ID>DATA_IN_7</ID>528 </input>
<output>
<ID>DATA_OUT_0</ID>537 </output>
<output>
<ID>DATA_OUT_1</ID>522 </output>
<output>
<ID>DATA_OUT_2</ID>523 </output>
<output>
<ID>DATA_OUT_3</ID>524 </output>
<output>
<ID>DATA_OUT_4</ID>525 </output>
<output>
<ID>DATA_OUT_5</ID>526 </output>
<output>
<ID>DATA_OUT_6</ID>527 </output>
<output>
<ID>DATA_OUT_7</ID>528 </output>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>write_enable</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_REGISTER8</type>
<position>65,-32.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>513 </input>
<input>
<ID>IN_2</ID>512 </input>
<input>
<ID>IN_3</ID>511 </input>
<input>
<ID>IN_4</ID>510 </input>
<input>
<ID>IN_5</ID>509 </input>
<input>
<ID>IN_6</ID>508 </input>
<input>
<ID>IN_7</ID>507 </input>
<output>
<ID>OUT_0</ID>516 </output>
<output>
<ID>OUT_1</ID>517 </output>
<input>
<ID>clear</ID>519 </input>
<input>
<ID>clock</ID>518 </input>
<input>
<ID>load</ID>515 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>352</ID>
<type>DD_KEYPAD_HEX</type>
<position>-24.5,-21</position>
<output>
<ID>OUT_0</ID>480 </output>
<output>
<ID>OUT_1</ID>481 </output>
<output>
<ID>OUT_2</ID>482 </output>
<output>
<ID>OUT_3</ID>483 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>353</ID>
<type>DD_KEYPAD_HEX</type>
<position>-24.5,-9</position>
<output>
<ID>OUT_0</ID>484 </output>
<output>
<ID>OUT_1</ID>485 </output>
<output>
<ID>OUT_2</ID>486 </output>
<output>
<ID>OUT_3</ID>487 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>354</ID>
<type>BB_CLOCK</type>
<position>-36,-46.5</position>
<output>
<ID>CLK</ID>539 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_TOGGLE</type>
<position>-7,4</position>
<output>
<ID>OUT_0</ID>503 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>-19.5,2</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>357</ID>
<type>AA_LABEL</type>
<position>-19.5,4.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>6,1.5</position>
<output>
<ID>OUT_0</ID>502 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_TOGGLE</type>
<position>-6,-43.5</position>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_LABEL</type>
<position>-11.5,-40.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>AA_TOGGLE</type>
<position>45,-25</position>
<output>
<ID>OUT_0</ID>504 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>-10,-7</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>6.5,-7</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_LABEL</type>
<position>27,-6</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>49,-22</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_TOGGLE</type>
<position>62,-24.5</position>
<output>
<ID>OUT_0</ID>515 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>367</ID>
<type>BE_ROM_8x8</type>
<position>80,-32</position>
<input>
<ID>ADDRESS_0</ID>516 </input>
<input>
<ID>ADDRESS_1</ID>517 </input>
<input>
<ID>ENABLE_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>368</ID>
<type>AA_TOGGLE</type>
<position>37,-12</position>
<output>
<ID>OUT_0</ID>520 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_TOGGLE</type>
<position>37,-15</position>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>43.5,-11.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>AA_LABEL</type>
<position>44,-14.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>41,-32</position>
<input>
<ID>ENABLE_0</ID>521 </input>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>522 </input>
<input>
<ID>IN_2</ID>523 </input>
<input>
<ID>IN_3</ID>524 </input>
<input>
<ID>IN_4</ID>525 </input>
<input>
<ID>IN_5</ID>526 </input>
<input>
<ID>IN_6</ID>527 </input>
<input>
<ID>IN_7</ID>528 </input>
<output>
<ID>OUT_0</ID>530 </output>
<output>
<ID>OUT_1</ID>531 </output>
<output>
<ID>OUT_2</ID>532 </output>
<output>
<ID>OUT_3</ID>533 </output>
<output>
<ID>OUT_4</ID>534 </output>
<output>
<ID>OUT_5</ID>529 </output>
<output>
<ID>OUT_6</ID>536 </output>
<output>
<ID>OUT_7</ID>535 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>373</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>20,-32</position>
<input>
<ID>ENABLE_0</ID>520 </input>
<output>
<ID>OUT_0</ID>537 </output>
<output>
<ID>OUT_1</ID>522 </output>
<output>
<ID>OUT_2</ID>523 </output>
<output>
<ID>OUT_3</ID>524 </output>
<output>
<ID>OUT_4</ID>525 </output>
<output>
<ID>OUT_5</ID>526 </output>
<output>
<ID>OUT_6</ID>527 </output>
<output>
<ID>OUT_7</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_LABEL</type>
<position>66.5,-24</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>375</ID>
<type>AA_TOGGLE</type>
<position>89,-32.5</position>
<output>
<ID>OUT_0</ID>538 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>376</ID>
<type>AA_LABEL</type>
<position>90.5,-29.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND2</type>
<position>-10,-28</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>542 </input>
<output>
<ID>OUT</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_AND2</type>
<position>-24.5,-45.5</position>
<input>
<ID>IN_0</ID>540 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AA_TOGGLE</type>
<position>-30,-42.5</position>
<output>
<ID>OUT_0</ID>540 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_TOGGLE</type>
<position>-39,-29</position>
<output>
<ID>OUT_0</ID>542 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>381</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>14,-87.5</position>
<input>
<ID>ENABLE_0</ID>563 </input>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>545 </input>
<input>
<ID>IN_10</ID>554 </input>
<input>
<ID>IN_11</ID>555 </input>
<input>
<ID>IN_12</ID>556 </input>
<input>
<ID>IN_13</ID>557 </input>
<input>
<ID>IN_14</ID>558 </input>
<input>
<ID>IN_15</ID>559 </input>
<input>
<ID>IN_2</ID>546 </input>
<input>
<ID>IN_3</ID>547 </input>
<input>
<ID>IN_4</ID>548 </input>
<input>
<ID>IN_5</ID>549 </input>
<input>
<ID>IN_6</ID>550 </input>
<input>
<ID>IN_7</ID>551 </input>
<input>
<ID>IN_8</ID>552 </input>
<input>
<ID>IN_9</ID>553 </input>
<output>
<ID>OUT_0</ID>581 </output>
<output>
<ID>OUT_1</ID>582 </output>
<output>
<ID>OUT_10</ID>591 </output>
<output>
<ID>OUT_11</ID>592 </output>
<output>
<ID>OUT_12</ID>593 </output>
<output>
<ID>OUT_13</ID>594 </output>
<output>
<ID>OUT_14</ID>595 </output>
<output>
<ID>OUT_15</ID>596 </output>
<output>
<ID>OUT_2</ID>583 </output>
<output>
<ID>OUT_3</ID>584 </output>
<output>
<ID>OUT_4</ID>585 </output>
<output>
<ID>OUT_5</ID>586 </output>
<output>
<ID>OUT_6</ID>587 </output>
<output>
<ID>OUT_7</ID>588 </output>
<output>
<ID>OUT_8</ID>589 </output>
<output>
<ID>OUT_9</ID>590 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>382</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>14,-110.5</position>
<input>
<ID>ENABLE_0</ID>562 </input>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>545 </input>
<input>
<ID>IN_10</ID>554 </input>
<input>
<ID>IN_11</ID>555 </input>
<input>
<ID>IN_12</ID>556 </input>
<input>
<ID>IN_13</ID>557 </input>
<input>
<ID>IN_14</ID>558 </input>
<input>
<ID>IN_15</ID>559 </input>
<input>
<ID>IN_2</ID>546 </input>
<input>
<ID>IN_3</ID>547 </input>
<input>
<ID>IN_4</ID>548 </input>
<input>
<ID>IN_5</ID>549 </input>
<input>
<ID>IN_6</ID>550 </input>
<input>
<ID>IN_7</ID>551 </input>
<input>
<ID>IN_8</ID>552 </input>
<input>
<ID>IN_9</ID>553 </input>
<output>
<ID>OUT_0</ID>565 </output>
<output>
<ID>OUT_1</ID>573 </output>
<output>
<ID>OUT_10</ID>570 </output>
<output>
<ID>OUT_11</ID>578 </output>
<output>
<ID>OUT_12</ID>571 </output>
<output>
<ID>OUT_13</ID>579 </output>
<output>
<ID>OUT_14</ID>572 </output>
<output>
<ID>OUT_15</ID>580 </output>
<output>
<ID>OUT_2</ID>566 </output>
<output>
<ID>OUT_3</ID>574 </output>
<output>
<ID>OUT_4</ID>567 </output>
<output>
<ID>OUT_5</ID>575 </output>
<output>
<ID>OUT_6</ID>568 </output>
<output>
<ID>OUT_7</ID>576 </output>
<output>
<ID>OUT_8</ID>569 </output>
<output>
<ID>OUT_9</ID>577 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_LABEL</type>
<position>-8.5,-74.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-81</position>
<output>
<ID>OUT_0</ID>553 </output>
<output>
<ID>OUT_1</ID>555 </output>
<output>
<ID>OUT_2</ID>557 </output>
<output>
<ID>OUT_3</ID>559 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>385</ID>
<type>DD_KEYPAD_HEX</type>
<position>-26,-105</position>
<output>
<ID>OUT_0</ID>552 </output>
<output>
<ID>OUT_1</ID>554 </output>
<output>
<ID>OUT_2</ID>556 </output>
<output>
<ID>OUT_3</ID>558 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-24,-14.5,-18</points>
<intersection>-24 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-18,-9,-18</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-24,-14.5,-24</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-22,-14.5,-17</points>
<intersection>-22 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-17,-9,-17</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-22,-14.5,-22</points>
<connection>
<GID>352</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-20,-14.5,-16</points>
<intersection>-20 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-16,-9,-16</points>
<connection>
<GID>347</GID>
<name>IN_2</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-20,-14.5,-20</points>
<connection>
<GID>352</GID>
<name>OUT_2</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-18,-14.5,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-15,-9,-15</points>
<connection>
<GID>347</GID>
<name>IN_3</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-18,-14.5,-18</points>
<connection>
<GID>352</GID>
<name>OUT_3</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-14,-14.5,-12</points>
<intersection>-14 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-14,-9,-14</points>
<connection>
<GID>347</GID>
<name>IN_4</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-12,-14.5,-12</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-13,-14.5,-10</points>
<intersection>-13 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-13,-9,-13</points>
<connection>
<GID>347</GID>
<name>IN_5</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-10,-14.5,-10</points>
<connection>
<GID>353</GID>
<name>OUT_1</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-12,-14.5,-8</points>
<intersection>-12 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,-12,-9,-12</points>
<connection>
<GID>347</GID>
<name>IN_6</name></connection>
<intersection>-14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-8,-14.5,-8</points>
<connection>
<GID>353</GID>
<name>OUT_2</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-11,-9,-11</points>
<connection>
<GID>347</GID>
<name>IN_7</name></connection>
<intersection>-19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19.5,-11,-19.5,-6</points>
<connection>
<GID>353</GID>
<name>OUT_3</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-11,8,-11</points>
<connection>
<GID>348</GID>
<name>IN_7</name></connection>
<connection>
<GID>347</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-12,8,-12</points>
<connection>
<GID>348</GID>
<name>IN_6</name></connection>
<connection>
<GID>347</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-13,8,-13</points>
<connection>
<GID>348</GID>
<name>IN_5</name></connection>
<connection>
<GID>347</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-14,8,-14</points>
<connection>
<GID>348</GID>
<name>IN_4</name></connection>
<connection>
<GID>347</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-15,8,-15</points>
<connection>
<GID>348</GID>
<name>IN_3</name></connection>
<connection>
<GID>347</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-16,8,-16</points>
<connection>
<GID>348</GID>
<name>IN_2</name></connection>
<connection>
<GID>347</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-17,8,-17</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<connection>
<GID>347</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-18,8,-18</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-11,22,-11</points>
<connection>
<GID>350</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>348</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-12,22,-12</points>
<connection>
<GID>350</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>348</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-13,22,-13</points>
<connection>
<GID>350</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>348</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-14,22,-14</points>
<connection>
<GID>350</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>348</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-15,22,-15</points>
<connection>
<GID>350</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>348</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-16,22,-16</points>
<connection>
<GID>350</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>348</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-9,11,1.5</points>
<connection>
<GID>348</GID>
<name>load</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,1.5,11,1.5</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-9,-5,4</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<connection>
<GID>347</GID>
<name>count_enable</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5,-8,-4,-8</points>
<intersection>-5 0</intersection>
<intersection>-4 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4,-9,-4,-8</points>
<connection>
<GID>347</GID>
<name>count_up</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>47,-25,48,-25</points>
<connection>
<GID>361</GID>
<name>OUT_0</name></connection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-26.5,48,-25</points>
<connection>
<GID>349</GID>
<name>load</name></connection>
<intersection>-25 2</intersection></vsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-17,22,-17</points>
<connection>
<GID>350</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>348</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-18,22,-18</points>
<connection>
<GID>350</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-28.5,61,-28.5</points>
<connection>
<GID>351</GID>
<name>IN_7</name></connection>
<connection>
<GID>349</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-29.5,61,-29.5</points>
<connection>
<GID>351</GID>
<name>IN_6</name></connection>
<connection>
<GID>349</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-30.5,61,-30.5</points>
<connection>
<GID>351</GID>
<name>IN_5</name></connection>
<connection>
<GID>349</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-31.5,61,-31.5</points>
<connection>
<GID>351</GID>
<name>IN_4</name></connection>
<connection>
<GID>349</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-32.5,61,-32.5</points>
<connection>
<GID>351</GID>
<name>IN_3</name></connection>
<connection>
<GID>349</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-33.5,61,-33.5</points>
<connection>
<GID>351</GID>
<name>IN_2</name></connection>
<connection>
<GID>349</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-34.5,61,-34.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<connection>
<GID>349</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-35.5,61,-35.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-26.5,64,-24.5</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<connection>
<GID>351</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-35.5,75,-35.5</points>
<connection>
<GID>367</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-34.5,75,-34.5</points>
<connection>
<GID>367</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>351</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-45.5,11,-20</points>
<connection>
<GID>348</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-45.5,64,-45.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>-19 6</intersection>
<intersection>11 0</intersection>
<intersection>48 5</intersection>
<intersection>64 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>64,-45.5,64,-37.5</points>
<connection>
<GID>351</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>48,-45.5,48,-37.5</points>
<connection>
<GID>349</GID>
<name>clock</name></connection>
<intersection>-45.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-19,-45.5,-19,-27</points>
<intersection>-45.5 1</intersection>
<intersection>-27 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-19,-27,-13,-27</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-19 6</intersection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-43.5,-4,-20</points>
<connection>
<GID>359</GID>
<name>OUT_0</name></connection>
<connection>
<GID>347</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-4,-43.5,66,-43.5</points>
<intersection>-4 0</intersection>
<intersection>13 3</intersection>
<intersection>50 7</intersection>
<intersection>66 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-43.5,13,-20</points>
<connection>
<GID>348</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>66,-43.5,66,-37.5</points>
<connection>
<GID>351</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>50,-43.5,50,-37.5</points>
<connection>
<GID>349</GID>
<name>clear</name></connection>
<intersection>-43.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-12,35,-12</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-27,33,-12</points>
<intersection>-27 4</intersection>
<intersection>-14 7</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-27,33,-27</points>
<connection>
<GID>373</GID>
<name>ENABLE_0</name></connection>
<intersection>33 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>32,-14,33,-14</points>
<connection>
<GID>350</GID>
<name>write_enable</name></connection>
<intersection>33 3</intersection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-15,35,-15</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>ENABLE_0</name></connection>
<intersection>35 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35,-27,35,-15</points>
<intersection>-27 6</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35,-27,41,-27</points>
<connection>
<GID>372</GID>
<name>ENABLE_0</name></connection>
<intersection>35 5</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-34.5,39,-34.5</points>
<connection>
<GID>373</GID>
<name>OUT_1</name></connection>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29.5,-34.5,29.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_1</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-33.5,39,-33.5</points>
<connection>
<GID>373</GID>
<name>OUT_2</name></connection>
<connection>
<GID>372</GID>
<name>IN_2</name></connection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,-33.5,28.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_2</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-32.5,39,-32.5</points>
<connection>
<GID>373</GID>
<name>OUT_3</name></connection>
<connection>
<GID>372</GID>
<name>IN_3</name></connection>
<intersection>27.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>27.5,-32.5,27.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_3</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-31.5,39,-31.5</points>
<connection>
<GID>373</GID>
<name>OUT_4</name></connection>
<connection>
<GID>372</GID>
<name>IN_4</name></connection>
<intersection>26.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26.5,-31.5,26.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_4</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-30.5,39,-30.5</points>
<connection>
<GID>373</GID>
<name>OUT_5</name></connection>
<connection>
<GID>372</GID>
<name>IN_5</name></connection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-30.5,25.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_5</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-29.5,39,-29.5</points>
<connection>
<GID>373</GID>
<name>OUT_6</name></connection>
<connection>
<GID>372</GID>
<name>IN_6</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-29.5,24.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_6</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-28.5,39,-28.5</points>
<connection>
<GID>373</GID>
<name>OUT_7</name></connection>
<connection>
<GID>372</GID>
<name>IN_7</name></connection>
<intersection>23.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-28.5,23.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_7</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-30.5,45,-30.5</points>
<connection>
<GID>372</GID>
<name>OUT_5</name></connection>
<connection>
<GID>349</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-35.5,45,-35.5</points>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection>
<connection>
<GID>349</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-34.5,45,-34.5</points>
<connection>
<GID>372</GID>
<name>OUT_1</name></connection>
<connection>
<GID>349</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-33.5,45,-33.5</points>
<connection>
<GID>372</GID>
<name>OUT_2</name></connection>
<connection>
<GID>349</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-32.5,45,-32.5</points>
<connection>
<GID>372</GID>
<name>OUT_3</name></connection>
<connection>
<GID>349</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-31.5,45,-31.5</points>
<connection>
<GID>372</GID>
<name>OUT_4</name></connection>
<connection>
<GID>349</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-28.5,45,-28.5</points>
<connection>
<GID>372</GID>
<name>OUT_7</name></connection>
<connection>
<GID>349</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-29.5,45,-29.5</points>
<connection>
<GID>372</GID>
<name>OUT_6</name></connection>
<connection>
<GID>349</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-35.5,39,-35.5</points>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-35.5,30.5,-21.5</points>
<connection>
<GID>350</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>350</GID>
<name>DATA_IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-32.5,87,-32.5</points>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection>
<connection>
<GID>367</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32,-46.5,-27.5,-46.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<connection>
<GID>354</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-44.5,-27.5,-42.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-42.5,-27.5,-42.5</points>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-28,-6,-20</points>
<connection>
<GID>347</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-28,-6,-28</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37,-29,-13,-29</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-34 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-34,-29,-34,-26.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-9,-6,-1</points>
<connection>
<GID>347</GID>
<name>load</name></connection>
<intersection>-1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-34,-20.5,-34,-1</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-34,-1,-6,-1</points>
<intersection>-34 1</intersection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-120,-4.5,-118</points>
<intersection>-120 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-118,12,-118</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-120,-4.5,-120</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-118,12,-95</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-118 1</intersection></vsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-117,-4.5,-94</points>
<intersection>-117 1</intersection>
<intersection>-96 2</intersection>
<intersection>-94 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-117,12,-117</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-96,-4.5,-96</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-94,12,-94</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-118,-4.5,-116</points>
<intersection>-118 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-116,12,-116</points>
<connection>
<GID>382</GID>
<name>IN_2</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-118,-4.5,-118</points>
<connection>
<GID>387</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-116,12,-93</points>
<connection>
<GID>381</GID>
<name>IN_2</name></connection>
<intersection>-116 1</intersection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-115,-4.5,-92</points>
<intersection>-115 1</intersection>
<intersection>-94 2</intersection>
<intersection>-92 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-115,12,-115</points>
<connection>
<GID>382</GID>
<name>IN_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-94,-4.5,-94</points>
<connection>
<GID>386</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-92,12,-92</points>
<connection>
<GID>381</GID>
<name>IN_3</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-116,-4.5,-114</points>
<intersection>-116 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-114,12,-114</points>
<connection>
<GID>382</GID>
<name>IN_4</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-116,-4.5,-116</points>
<connection>
<GID>387</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-114,12,-91</points>
<connection>
<GID>381</GID>
<name>IN_4</name></connection>
<intersection>-114 1</intersection></vsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-113,-4.5,-90</points>
<intersection>-113 1</intersection>
<intersection>-92 2</intersection>
<intersection>-90 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-113,12,-113</points>
<connection>
<GID>382</GID>
<name>IN_5</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-92,-4.5,-92</points>
<connection>
<GID>386</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-4.5,-90,12,-90</points>
<connection>
<GID>381</GID>
<name>IN_5</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-114,-4.5,-112</points>
<intersection>-114 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-112,12,-112</points>
<connection>
<GID>382</GID>
<name>IN_6</name></connection>
<intersection>-4.5 0</intersection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-114,-4.5,-114</points>
<connection>
<GID>387</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-112,12,-89</points>
<connection>
<GID>381</GID>
<name>IN_6</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-111,-4.5,-88</points>
<intersection>-111 1</intersection>
<intersection>-90 2</intersection>
<intersection>-88 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-111,12,-111</points>
<connection>
<GID>382</GID>
<name>IN_7</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-90,-4.5,-90</points>
<connection>
<GID>386</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-88,12,-88</points>
<connection>
<GID>381</GID>
<name>IN_7</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-110,-4.5,-87</points>
<intersection>-110 1</intersection>
<intersection>-108 2</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-110,12,-110</points>
<connection>
<GID>382</GID>
<name>IN_8</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-108,-4.5,-108</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-87,12,-87</points>
<connection>
<GID>381</GID>
<name>IN_8</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-109,-4.5,-84</points>
<intersection>-109 1</intersection>
<intersection>-86 4</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-109,12,-109</points>
<connection>
<GID>382</GID>
<name>IN_9</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-84,-4.5,-84</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-86,12,-86</points>
<connection>
<GID>381</GID>
<name>IN_9</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-108,-4.5,-85</points>
<intersection>-108 1</intersection>
<intersection>-106 2</intersection>
<intersection>-85 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-108,12,-108</points>
<connection>
<GID>382</GID>
<name>IN_10</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-106,-4.5,-106</points>
<connection>
<GID>385</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-85,12,-85</points>
<connection>
<GID>381</GID>
<name>IN_10</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-107,-4.5,-82</points>
<intersection>-107 1</intersection>
<intersection>-84 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-107,12,-107</points>
<connection>
<GID>382</GID>
<name>IN_11</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-82,-4.5,-82</points>
<connection>
<GID>384</GID>
<name>OUT_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-84,12,-84</points>
<connection>
<GID>381</GID>
<name>IN_11</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-106,-4.5,-83</points>
<intersection>-106 1</intersection>
<intersection>-104 2</intersection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-106,12,-106</points>
<connection>
<GID>382</GID>
<name>IN_12</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-104,-4.5,-104</points>
<connection>
<GID>385</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-83,12,-83</points>
<connection>
<GID>381</GID>
<name>IN_12</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-105,-4.5,-80</points>
<intersection>-105 1</intersection>
<intersection>-82 3</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-105,12,-105</points>
<connection>
<GID>382</GID>
<name>IN_13</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-80,-4.5,-80</points>
<connection>
<GID>384</GID>
<name>OUT_2</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-82,12,-82</points>
<connection>
<GID>381</GID>
<name>IN_13</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-104,-4.5,-81</points>
<intersection>-104 1</intersection>
<intersection>-102 2</intersection>
<intersection>-81 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-104,12,-104</points>
<connection>
<GID>382</GID>
<name>IN_14</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-102,-4.5,-102</points>
<connection>
<GID>385</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-81,12,-81</points>
<connection>
<GID>381</GID>
<name>IN_14</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-103,-4.5,-78</points>
<intersection>-103 1</intersection>
<intersection>-80 3</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-103,12,-103</points>
<connection>
<GID>382</GID>
<name>IN_15</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-78,-4.5,-78</points>
<connection>
<GID>384</GID>
<name>OUT_3</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-80,12,-80</points>
<connection>
<GID>381</GID>
<name>IN_15</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-69.5,2.5,-69.5</points>
<connection>
<GID>392</GID>
<name>ENABLE</name></connection>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-64,54,-64</points>
<intersection>-2 8</intersection>
<intersection>54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>54,-115.5,54,-64</points>
<intersection>-115.5 18</intersection>
<intersection>-110.5 19</intersection>
<intersection>-105.5 20</intersection>
<intersection>-100.5 21</intersection>
<intersection>-95.5 22</intersection>
<intersection>-90.5 23</intersection>
<intersection>-85.5 24</intersection>
<intersection>-80.5 25</intersection>
<intersection>-64 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-2,-72.5,-2,-64</points>
<intersection>-72.5 10</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-2,-72.5,2.5,-72.5</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-2 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>54,-115.5,57,-115.5</points>
<connection>
<GID>420</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>54,-110.5,57,-110.5</points>
<connection>
<GID>419</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>54,-105.5,57,-105.5</points>
<connection>
<GID>418</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>54,-100.5,57,-100.5</points>
<connection>
<GID>417</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>54,-95.5,57,-95.5</points>
<connection>
<GID>416</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>54,-90.5,57,-90.5</points>
<connection>
<GID>415</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>54,-85.5,57,-85.5</points>
<connection>
<GID>414</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>54,-80.5,57,-80.5</points>
<connection>
<GID>413</GID>
<name>SEL_0</name></connection>
<intersection>54 7</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-101.5,9.5,-72.5</points>
<intersection>-101.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-72.5,9.5,-72.5</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-101.5,14,-101.5</points>
<connection>
<GID>382</GID>
<name>ENABLE_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-78.5,14,-71.5</points>
<connection>
<GID>381</GID>
<name>ENABLE_0</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-71.5,14,-71.5</points>
<connection>
<GID>392</GID>
<name>OUT_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-114.5,30.5,-114.5</points>
<connection>
<GID>397</GID>
<name>carry_out</name></connection>
<connection>
<GID>398</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-118,17.5,-101.5</points>
<intersection>-118 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-101.5,27.5,-101.5</points>
<connection>
<GID>397</GID>
<name>IN_B_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-118,17.5,-118</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-116,18,-102.5</points>
<intersection>-116 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-102.5,27.5,-102.5</points>
<connection>
<GID>397</GID>
<name>IN_B_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-116,18,-116</points>
<connection>
<GID>382</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-114,18.5,-103.5</points>
<intersection>-114 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-103.5,27.5,-103.5</points>
<connection>
<GID>397</GID>
<name>IN_B_2</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-114,18.5,-114</points>
<connection>
<GID>382</GID>
<name>OUT_4</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-112,19,-104.5</points>
<intersection>-112 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-104.5,27.5,-104.5</points>
<connection>
<GID>397</GID>
<name>IN_B_3</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-112,19,-112</points>
<connection>
<GID>382</GID>
<name>OUT_6</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-117.5,21,-110</points>
<intersection>-117.5 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-117.5,27.5,-117.5</points>
<connection>
<GID>398</GID>
<name>IN_B_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-110,21,-110</points>
<connection>
<GID>382</GID>
<name>OUT_8</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-118.5,20.5,-108</points>
<intersection>-118.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-118.5,27.5,-118.5</points>
<connection>
<GID>398</GID>
<name>IN_B_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-108,20.5,-108</points>
<connection>
<GID>382</GID>
<name>OUT_10</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-119.5,20,-106</points>
<intersection>-119.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-119.5,27.5,-119.5</points>
<connection>
<GID>398</GID>
<name>IN_B_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-106,20,-106</points>
<connection>
<GID>382</GID>
<name>OUT_12</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-120.5,19.5,-104</points>
<intersection>-120.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-120.5,27.5,-120.5</points>
<connection>
<GID>398</GID>
<name>IN_B_3</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-104,19.5,-104</points>
<connection>
<GID>382</GID>
<name>OUT_14</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-117,21.5,-108.5</points>
<intersection>-117 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-108.5,27.5,-108.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-117,21.5,-117</points>
<connection>
<GID>382</GID>
<name>OUT_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-115,21.5,-109.5</points>
<intersection>-115 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-109.5,27.5,-109.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-115,21.5,-115</points>
<connection>
<GID>382</GID>
<name>OUT_3</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-113,21.5,-110.5</points>
<intersection>-113 2</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-110.5,27.5,-110.5</points>
<connection>
<GID>397</GID>
<name>IN_2</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-113,21.5,-113</points>
<connection>
<GID>382</GID>
<name>OUT_5</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-111.5,21.5,-111</points>
<intersection>-111.5 1</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-111.5,27.5,-111.5</points>
<connection>
<GID>397</GID>
<name>IN_3</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-111,21.5,-111</points>
<connection>
<GID>382</GID>
<name>OUT_7</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-124.5,23.5,-109</points>
<intersection>-124.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-124.5,27.5,-124.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-109,23.5,-109</points>
<connection>
<GID>382</GID>
<name>OUT_9</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-125.5,23,-107</points>
<intersection>-125.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-125.5,27.5,-125.5</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-107,23,-107</points>
<connection>
<GID>382</GID>
<name>OUT_11</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-126.5,22.5,-105</points>
<intersection>-126.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-126.5,27.5,-126.5</points>
<connection>
<GID>398</GID>
<name>IN_2</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-105,22.5,-105</points>
<connection>
<GID>382</GID>
<name>OUT_13</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-127.5,22,-103</points>
<intersection>-127.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-127.5,27.5,-127.5</points>
<connection>
<GID>398</GID>
<name>IN_3</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-103,22,-103</points>
<connection>
<GID>382</GID>
<name>OUT_15</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-97,17,-95</points>
<intersection>-97 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-97,24,-97</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-95,17,-95</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-95,24,-95</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-95,16,-94</points>
<connection>
<GID>381</GID>
<name>OUT_1</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-93.5,19.5,-93</points>
<intersection>-93.5 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-93.5,29,-93.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-93,19.5,-93</points>
<connection>
<GID>381</GID>
<name>OUT_2</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-91.5,29,-91.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-92,16,-91.5</points>
<connection>
<GID>381</GID>
<name>OUT_3</name></connection>
<intersection>-91.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-90,24,-90</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-91,16,-90</points>
<connection>
<GID>381</GID>
<name>OUT_4</name></connection>
<intersection>-90 1</intersection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-90,17,-88</points>
<intersection>-90 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-88,24,-88</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-90,17,-90</points>
<connection>
<GID>381</GID>
<name>OUT_5</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-89,18,-86.5</points>
<intersection>-89 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-86.5,29,-86.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-89,18,-89</points>
<connection>
<GID>381</GID>
<name>OUT_6</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-88,17.5,-84.5</points>
<intersection>-88 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-84.5,29,-84.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-88,17.5,-88</points>
<connection>
<GID>381</GID>
<name>OUT_7</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-87,17,-83</points>
<intersection>-87 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-83,24,-83</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-87,17,-87</points>
<connection>
<GID>381</GID>
<name>OUT_8</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-86,17,-81</points>
<intersection>-86 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-81,24,-81</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-86,17,-86</points>
<connection>
<GID>381</GID>
<name>OUT_9</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-85,17.5,-79.5</points>
<intersection>-85 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-79.5,29,-79.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-85,17.5,-85</points>
<connection>
<GID>381</GID>
<name>OUT_10</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-84,17.5,-77.5</points>
<intersection>-84 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-77.5,29,-77.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-84,17.5,-84</points>
<connection>
<GID>381</GID>
<name>OUT_11</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-83,17,-76</points>
<intersection>-83 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-76,24,-76</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-83,17,-83</points>
<connection>
<GID>381</GID>
<name>OUT_12</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-82,17,-74</points>
<intersection>-82 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-74,24,-74</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-82,17,-82</points>
<connection>
<GID>381</GID>
<name>OUT_13</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-81,16.5,-72.5</points>
<intersection>-81 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-72.5,29,-72.5</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-81,16.5,-81</points>
<connection>
<GID>381</GID>
<name>OUT_14</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-80,16,-70.5</points>
<connection>
<GID>381</GID>
<name>OUT_15</name></connection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-70.5,29,-70.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-119,45,-105</points>
<intersection>-119 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-119,55,-119</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-105,45,-105</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-114,45,-106</points>
<intersection>-114 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-114,55,-114</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-106,45,-106</points>
<connection>
<GID>397</GID>
<name>OUT_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-109,45,-107</points>
<intersection>-109 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-109,55,-109</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-107,45,-107</points>
<connection>
<GID>397</GID>
<name>OUT_2</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-108,45,-104</points>
<intersection>-108 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-104,55,-104</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-108,45,-108</points>
<connection>
<GID>397</GID>
<name>OUT_3</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-121,45,-99</points>
<intersection>-121 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-99,55,-99</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-121,45,-121</points>
<connection>
<GID>398</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-122,45,-94</points>
<intersection>-122 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-94,55,-94</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-122,45,-122</points>
<connection>
<GID>398</GID>
<name>OUT_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-123,45,-89</points>
<intersection>-123 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-89,55,-89</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-123,45,-123</points>
<connection>
<GID>398</GID>
<name>OUT_2</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-124,45,-84</points>
<intersection>-124 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-84,55,-84</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-124,45,-124</points>
<connection>
<GID>398</GID>
<name>OUT_3</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-117,42.5,-96</points>
<intersection>-117 1</intersection>
<intersection>-96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-117,55,-117</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-96,42.5,-96</points>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-112,45,-92.5</points>
<intersection>-112 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-92.5,45,-92.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-112,55,-112</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-107,42.5,-89</points>
<intersection>-107 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-89,42.5,-89</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-107,55,-107</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-102,45,-85.5</points>
<intersection>-102 2</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-85.5,45,-85.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-102,55,-102</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-97,42.5,-82</points>
<intersection>-97 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-82,42.5,-82</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-97,55,-97</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-92,45,-78.5</points>
<intersection>-92 2</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-78.5,45,-78.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-92,55,-92</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-87,42.5,-75</points>
<intersection>-87 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-75,42.5,-75</points>
<connection>
<GID>411</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-87,55,-87</points>
<connection>
<GID>414</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-82,45,-71.5</points>
<intersection>-82 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-71.5,45,-71.5</points>
<connection>
<GID>412</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-82,55,-82</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-118,66.5,-103</points>
<intersection>-118 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-103,74.5,-103</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection>
<intersection>67.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-118,66.5,-118</points>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>67.5,-108.5,67.5,-103</points>
<intersection>-108.5 8</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>67.5,-108.5,88.5,-108.5</points>
<intersection>67.5 7</intersection>
<intersection>88.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>88.5,-109,88.5,-108.5</points>
<connection>
<GID>431</GID>
<name>N_in2</name></connection>
<intersection>-108.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-113,66.5,-102</points>
<intersection>-113 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-102,74.5,-102</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>66.5 0</intersection>
<intersection>68 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-113,66.5,-113</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>68,-108,68,-102</points>
<intersection>-108 8</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68,-108,86,-108</points>
<intersection>68 7</intersection>
<intersection>86 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>86,-109,86,-108</points>
<connection>
<GID>430</GID>
<name>N_in2</name></connection>
<intersection>-108 8</intersection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-108,66.5,-101</points>
<intersection>-108 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-101,74.5,-101</points>
<connection>
<GID>421</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection>
<intersection>68.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-108,66.5,-108</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>68.5,-107.5,68.5,-101</points>
<intersection>-107.5 8</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-107.5,83.5,-107.5</points>
<intersection>68.5 7</intersection>
<intersection>83.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>83.5,-109,83.5,-107.5</points>
<connection>
<GID>429</GID>
<name>N_in2</name></connection>
<intersection>-107.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-103,66.5,-100</points>
<intersection>-103 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-100,74.5,-100</points>
<connection>
<GID>421</GID>
<name>IN_3</name></connection>
<intersection>66.5 0</intersection>
<intersection>69 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-103,66.5,-103</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>69,-107,69,-100</points>
<intersection>-107 9</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>69,-107,81,-107</points>
<intersection>69 8</intersection>
<intersection>81 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>81,-109,81,-107</points>
<connection>
<GID>428</GID>
<name>N_in2</name></connection>
<intersection>-107 9</intersection></vsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-99,66.5,-98</points>
<intersection>-99 1</intersection>
<intersection>-98 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-99,74.5,-99</points>
<connection>
<GID>421</GID>
<name>IN_4</name></connection>
<intersection>66.5 0</intersection>
<intersection>69.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-98,66.5,-98</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>69.5,-106.5,69.5,-99</points>
<intersection>-106.5 9</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>69.5,-106.5,78.5,-106.5</points>
<intersection>69.5 8</intersection>
<intersection>78.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>78.5,-109,78.5,-106.5</points>
<connection>
<GID>427</GID>
<name>N_in2</name></connection>
<intersection>-106.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-98,66.5,-93</points>
<intersection>-98 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-98,74.5,-98</points>
<connection>
<GID>421</GID>
<name>IN_5</name></connection>
<intersection>66.5 0</intersection>
<intersection>70 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-93,66.5,-93</points>
<connection>
<GID>415</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70,-106,70,-98</points>
<intersection>-106 8</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>70,-106,76,-106</points>
<intersection>70 7</intersection>
<intersection>76 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>76,-109,76,-106</points>
<connection>
<GID>426</GID>
<name>N_in2</name></connection>
<intersection>-106 8</intersection></vsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-97,66.5,-88</points>
<intersection>-97 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-97,74.5,-97</points>
<connection>
<GID>421</GID>
<name>IN_6</name></connection>
<intersection>66.5 0</intersection>
<intersection>70.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-88,66.5,-88</points>
<connection>
<GID>414</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70.5,-105.5,70.5,-97</points>
<intersection>-105.5 8</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>70.5,-105.5,73.5,-105.5</points>
<intersection>70.5 7</intersection>
<intersection>73.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>73.5,-109,73.5,-105.5</points>
<connection>
<GID>425</GID>
<name>N_in2</name></connection>
<intersection>-105.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-96,66.5,-83</points>
<intersection>-96 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-83,66.5,-83</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-96,74.5,-96</points>
<connection>
<GID>421</GID>
<name>IN_7</name></connection>
<intersection>66.5 0</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71,-109,71,-96</points>
<connection>
<GID>424</GID>
<name>N_in2</name></connection>
<intersection>-96 2</intersection></vsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-44,172,-44</points>
<connection>
<GID>479</GID>
<name>OUT_7</name></connection>
<intersection>172 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>172,-44,172,-34</points>
<intersection>-44 1</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>172,-34,185,-34</points>
<connection>
<GID>461</GID>
<name>IN_3</name></connection>
<connection>
<GID>444</GID>
<name>IN_3</name></connection>
<intersection>172 4</intersection>
<intersection>183.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>183.5,-40,183.5,-34</points>
<intersection>-40 8</intersection>
<intersection>-34 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>183.5,-40,185,-40</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>183.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-45,185,-45</points>
<connection>
<GID>479</GID>
<name>OUT_6</name></connection>
<connection>
<GID>462</GID>
<name>IN_3</name></connection>
<connection>
<GID>445</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-56,171,-46</points>
<intersection>-56 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-56,185,-56</points>
<connection>
<GID>463</GID>
<name>IN_3</name></connection>
<connection>
<GID>446</GID>
<name>IN_3</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-46,171,-46</points>
<connection>
<GID>479</GID>
<name>OUT_5</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-65.5,170.5,-47</points>
<intersection>-65.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-65.5,185,-65.5</points>
<connection>
<GID>464</GID>
<name>IN_3</name></connection>
<connection>
<GID>447</GID>
<name>IN_3</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-47,170.5,-47</points>
<connection>
<GID>479</GID>
<name>OUT_4</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-76.5,170,-48</points>
<intersection>-76.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-76.5,185,-76.5</points>
<connection>
<GID>465</GID>
<name>IN_3</name></connection>
<connection>
<GID>448</GID>
<name>IN_3</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-48,170,-48</points>
<connection>
<GID>479</GID>
<name>OUT_3</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-87.5,169.5,-49</points>
<intersection>-87.5 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-87.5,185,-87.5</points>
<connection>
<GID>466</GID>
<name>IN_3</name></connection>
<connection>
<GID>449</GID>
<name>IN_3</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-49,169.5,-49</points>
<connection>
<GID>479</GID>
<name>OUT_2</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-98,169,-50</points>
<intersection>-98 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169,-98,185,-98</points>
<connection>
<GID>467</GID>
<name>IN_3</name></connection>
<connection>
<GID>450</GID>
<name>IN_3</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-50,169,-50</points>
<connection>
<GID>479</GID>
<name>OUT_1</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-109,168.5,-51</points>
<intersection>-109 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-51,168.5,-51</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-109,185,-109</points>
<connection>
<GID>468</GID>
<name>IN_3</name></connection>
<connection>
<GID>451</GID>
<name>IN_3</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-57,167.5,-36</points>
<intersection>-57 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-36,185,-36</points>
<connection>
<GID>461</GID>
<name>IN_2</name></connection>
<connection>
<GID>444</GID>
<name>IN_2</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-57,167.5,-57</points>
<connection>
<GID>480</GID>
<name>OUT_7</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-58,167,-47</points>
<intersection>-58 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-47,185,-47</points>
<connection>
<GID>462</GID>
<name>IN_2</name></connection>
<connection>
<GID>445</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-58,167,-58</points>
<connection>
<GID>480</GID>
<name>OUT_6</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-59,172.5,-59</points>
<connection>
<GID>480</GID>
<name>OUT_5</name></connection>
<intersection>172.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>172.5,-59,172.5,-58</points>
<connection>
<GID>446</GID>
<name>IN_2</name></connection>
<intersection>-59 1</intersection>
<intersection>-58 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-58,185,-58</points>
<connection>
<GID>463</GID>
<name>IN_2</name></connection>
<intersection>172.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-67.5,166.5,-60</points>
<intersection>-67.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-67.5,185,-67.5</points>
<connection>
<GID>464</GID>
<name>IN_2</name></connection>
<connection>
<GID>447</GID>
<name>IN_2</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-60,166.5,-60</points>
<connection>
<GID>480</GID>
<name>OUT_4</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-78.5,166,-61</points>
<intersection>-78.5 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-78.5,185,-78.5</points>
<connection>
<GID>465</GID>
<name>IN_2</name></connection>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-61,166,-61</points>
<connection>
<GID>480</GID>
<name>OUT_3</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-89.5,165.5,-62</points>
<intersection>-89.5 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165.5,-89.5,185,-89.5</points>
<connection>
<GID>466</GID>
<name>IN_2</name></connection>
<connection>
<GID>449</GID>
<name>IN_2</name></connection>
<intersection>165.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-62,165.5,-62</points>
<connection>
<GID>480</GID>
<name>OUT_2</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165,-100,165,-63</points>
<intersection>-100 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-63,165,-63</points>
<connection>
<GID>480</GID>
<name>OUT_1</name></connection>
<intersection>165 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-100,185,-100</points>
<connection>
<GID>467</GID>
<name>IN_2</name></connection>
<connection>
<GID>450</GID>
<name>IN_2</name></connection>
<intersection>165 0</intersection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-111,168,-64</points>
<intersection>-111 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-111,185,-111</points>
<connection>
<GID>468</GID>
<name>IN_2</name></connection>
<connection>
<GID>451</GID>
<name>IN_2</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-64,168,-64</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-70.5,163.5,-38</points>
<intersection>-70.5 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-38,185,-38</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-70.5,163.5,-70.5</points>
<connection>
<GID>442</GID>
<name>OUT_7</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-71.5,163,-49</points>
<intersection>-71.5 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-49,185,-49</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-71.5,163,-71.5</points>
<connection>
<GID>442</GID>
<name>OUT_6</name></connection>
<intersection>163 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-72.5,162.5,-60</points>
<intersection>-72.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-60,185,-60</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>162.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-72.5,162.5,-72.5</points>
<connection>
<GID>442</GID>
<name>OUT_5</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-73.5,162,-69.5</points>
<intersection>-73.5 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-69.5,185,-69.5</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-73.5,162,-73.5</points>
<connection>
<GID>442</GID>
<name>OUT_4</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-80.5,161.5,-74.5</points>
<intersection>-80.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-80.5,185,-80.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>161.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-74.5,161.5,-74.5</points>
<connection>
<GID>442</GID>
<name>OUT_3</name></connection>
<intersection>161.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-91.5,161,-75.5</points>
<intersection>-91.5 1</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-91.5,185,-91.5</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-75.5,161,-75.5</points>
<connection>
<GID>442</GID>
<name>OUT_2</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-102,160.5,-76.5</points>
<intersection>-102 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-102,185,-102</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-76.5,160.5,-76.5</points>
<connection>
<GID>442</GID>
<name>OUT_1</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-113,160,-77.5</points>
<intersection>-113 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-77.5,160,-77.5</points>
<connection>
<GID>442</GID>
<name>OUT_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-113,185,-113</points>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<connection>
<GID>451</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-83.5,159,-40</points>
<intersection>-83.5 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159,-40,172.5,-40</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-83.5,159,-83.5</points>
<connection>
<GID>443</GID>
<name>OUT_7</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-84.5,158.5,-51</points>
<intersection>-84.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,-51,185,-51</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-84.5,158.5,-84.5</points>
<connection>
<GID>443</GID>
<name>OUT_6</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-85.5,158,-62</points>
<intersection>-85.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,-62,185,-62</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-85.5,158,-85.5</points>
<connection>
<GID>443</GID>
<name>OUT_5</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-71.5,185,-71.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>154 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>154,-86.5,154,-71.5</points>
<connection>
<GID>443</GID>
<name>OUT_4</name></connection>
<intersection>-71.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-87.5,157,-82.5</points>
<intersection>-87.5 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-82.5,185,-82.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-87.5,157,-87.5</points>
<connection>
<GID>443</GID>
<name>OUT_3</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-93.5,156.5,-88.5</points>
<intersection>-93.5 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-93.5,185,-93.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-88.5,156.5,-88.5</points>
<connection>
<GID>443</GID>
<name>OUT_2</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-104,156,-89.5</points>
<intersection>-104 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-104,185,-104</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-89.5,156,-89.5</points>
<connection>
<GID>443</GID>
<name>OUT_1</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-65.5,197,-37</points>
<intersection>-65.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-37,197,-37</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-65.5,202.5,-65.5</points>
<connection>
<GID>452</GID>
<name>IN_7</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-66.5,197,-48</points>
<intersection>-66.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-48,197,-48</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-66.5,202.5,-66.5</points>
<connection>
<GID>452</GID>
<name>IN_6</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-67.5,197,-59</points>
<intersection>-67.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-59,197,-59</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-67.5,202.5,-67.5</points>
<connection>
<GID>452</GID>
<name>IN_5</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>178.5,-68.5,202.5,-68.5</points>
<connection>
<GID>452</GID>
<name>IN_4</name></connection>
<connection>
<GID>447</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-79.5,197,-69.5</points>
<intersection>-79.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-79.5,197,-79.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-69.5,202.5,-69.5</points>
<connection>
<GID>452</GID>
<name>IN_3</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-90.5,197,-70.5</points>
<intersection>-90.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-90.5,197,-90.5</points>
<connection>
<GID>449</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-70.5,202.5,-70.5</points>
<connection>
<GID>452</GID>
<name>IN_2</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-101,197,-71.5</points>
<intersection>-101 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-101,197,-101</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-71.5,202.5,-71.5</points>
<connection>
<GID>452</GID>
<name>IN_1</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-112,197,-72.5</points>
<intersection>-112 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-72.5,202.5,-72.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-112,197,-112</points>
<connection>
<GID>451</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-115,155.5,-90.5</points>
<intersection>-115 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-115,185,-115</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-90.5,155.5,-90.5</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-96,145.5,-53</points>
<intersection>-96 10</intersection>
<intersection>-92.5 8</intersection>
<intersection>-79.5 7</intersection>
<intersection>-66 6</intersection>
<intersection>-53 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>145.5,-53,149,-53</points>
<connection>
<GID>479</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>145.5,-66,149,-66</points>
<connection>
<GID>480</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>145.5,-79.5,149,-79.5</points>
<connection>
<GID>442</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>145.5,-92.5,149,-92.5</points>
<connection>
<GID>443</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>142.5,-96,145.5,-96</points>
<connection>
<GID>454</GID>
<name>CLK</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-107,176.5,-29</points>
<connection>
<GID>451</GID>
<name>SEL_0</name></connection>
<connection>
<GID>450</GID>
<name>SEL_0</name></connection>
<connection>
<GID>449</GID>
<name>SEL_0</name></connection>
<connection>
<GID>448</GID>
<name>SEL_0</name></connection>
<connection>
<GID>447</GID>
<name>SEL_0</name></connection>
<connection>
<GID>446</GID>
<name>SEL_0</name></connection>
<connection>
<GID>445</GID>
<name>SEL_0</name></connection>
<connection>
<GID>444</GID>
<name>SEL_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-29,176.5,-29</points>
<intersection>123 2</intersection>
<intersection>176.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>123,-55,123,-29</points>
<intersection>-55 3</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-55,123,-55</points>
<connection>
<GID>453</GID>
<name>OUT_0</name></connection>
<intersection>123 2</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-107,175.5,-29.5</points>
<connection>
<GID>451</GID>
<name>SEL_1</name></connection>
<connection>
<GID>450</GID>
<name>SEL_1</name></connection>
<connection>
<GID>449</GID>
<name>SEL_1</name></connection>
<connection>
<GID>448</GID>
<name>SEL_1</name></connection>
<connection>
<GID>447</GID>
<name>SEL_1</name></connection>
<connection>
<GID>446</GID>
<name>SEL_1</name></connection>
<connection>
<GID>445</GID>
<name>SEL_1</name></connection>
<connection>
<GID>444</GID>
<name>SEL_1</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-29.5,175.5,-29.5</points>
<intersection>122.5 2</intersection>
<intersection>175.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>122.5,-53,122.5,-29.5</points>
<intersection>-53 3</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-53,122.5,-53</points>
<connection>
<GID>453</GID>
<name>OUT_1</name></connection>
<intersection>122.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-76.5,191.5,-37</points>
<intersection>-76.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-37,191.5,-37</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-76.5,202.5,-76.5</points>
<connection>
<GID>469</GID>
<name>IN_7</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-77.5,191.5,-48</points>
<intersection>-77.5 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-48,191.5,-48</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-77.5,202.5,-77.5</points>
<connection>
<GID>469</GID>
<name>IN_6</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-78.5,191.5,-59</points>
<intersection>-78.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-59,191.5,-59</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-78.5,202.5,-78.5</points>
<connection>
<GID>469</GID>
<name>IN_5</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-79.5,191.5,-68.5</points>
<intersection>-79.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-68.5,191.5,-68.5</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-79.5,202.5,-79.5</points>
<connection>
<GID>469</GID>
<name>IN_4</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-80.5,202.5,-80.5</points>
<connection>
<GID>469</GID>
<name>IN_3</name></connection>
<intersection>191.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>191.5,-80.5,191.5,-79.5</points>
<intersection>-80.5 1</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>191,-79.5,191.5,-79.5</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>191.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-90.5,191.5,-81.5</points>
<intersection>-90.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-90.5,191.5,-90.5</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-81.5,202.5,-81.5</points>
<connection>
<GID>469</GID>
<name>IN_2</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-101,191.5,-82.5</points>
<intersection>-101 1</intersection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-101,191.5,-101</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-82.5,202.5,-82.5</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-112,191.5,-83.5</points>
<intersection>-112 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-83.5,202.5,-83.5</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-112,191.5,-112</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-107,189,-30.5</points>
<connection>
<GID>468</GID>
<name>SEL_0</name></connection>
<connection>
<GID>467</GID>
<name>SEL_0</name></connection>
<connection>
<GID>466</GID>
<name>SEL_0</name></connection>
<connection>
<GID>465</GID>
<name>SEL_0</name></connection>
<connection>
<GID>464</GID>
<name>SEL_0</name></connection>
<connection>
<GID>463</GID>
<name>SEL_0</name></connection>
<connection>
<GID>462</GID>
<name>SEL_0</name></connection>
<connection>
<GID>461</GID>
<name>SEL_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-30.5,189,-30.5</points>
<intersection>124 2</intersection>
<intersection>189 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124,-69,124,-30.5</points>
<intersection>-69 3</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122,-69,124,-69</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>124 2</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-107,188,-30</points>
<connection>
<GID>468</GID>
<name>SEL_1</name></connection>
<connection>
<GID>467</GID>
<name>SEL_1</name></connection>
<connection>
<GID>466</GID>
<name>SEL_1</name></connection>
<connection>
<GID>465</GID>
<name>SEL_1</name></connection>
<connection>
<GID>464</GID>
<name>SEL_1</name></connection>
<connection>
<GID>463</GID>
<name>SEL_1</name></connection>
<connection>
<GID>462</GID>
<name>SEL_1</name></connection>
<connection>
<GID>461</GID>
<name>SEL_1</name></connection>
<intersection>-30 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>123.5,-30,188,-30</points>
<intersection>123.5 16</intersection>
<intersection>188 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>123.5,-67,123.5,-30</points>
<intersection>-67 18</intersection>
<intersection>-30 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>122,-67,123.5,-67</points>
<connection>
<GID>460</GID>
<name>OUT_1</name></connection>
<intersection>123.5 16</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-83.5,144.5,-44</points>
<intersection>-83.5 6</intersection>
<intersection>-70.5 3</intersection>
<intersection>-62.5 4</intersection>
<intersection>-57 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-44,146,-44</points>
<connection>
<GID>479</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-57,146,-57</points>
<connection>
<GID>480</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144.5,-70.5,146,-70.5</points>
<connection>
<GID>442</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>138,-62.5,144.5,-62.5</points>
<connection>
<GID>471</GID>
<name>OUT_3</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>144.5,-83.5,146,-83.5</points>
<connection>
<GID>443</GID>
<name>IN_7</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-84.5,144,-45</points>
<intersection>-84.5 6</intersection>
<intersection>-71.5 5</intersection>
<intersection>-64.5 2</intersection>
<intersection>-58 3</intersection>
<intersection>-45 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-64.5,144,-64.5</points>
<connection>
<GID>471</GID>
<name>OUT_2</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144,-58,146,-58</points>
<connection>
<GID>480</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>144,-45,146,-45</points>
<connection>
<GID>479</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>144,-71.5,146,-71.5</points>
<connection>
<GID>442</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>144,-84.5,146,-84.5</points>
<connection>
<GID>443</GID>
<name>IN_6</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-85.5,143.5,-46</points>
<intersection>-85.5 6</intersection>
<intersection>-72.5 3</intersection>
<intersection>-66.5 2</intersection>
<intersection>-59 4</intersection>
<intersection>-46 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-66.5,143.5,-66.5</points>
<connection>
<GID>471</GID>
<name>OUT_1</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>143.5,-72.5,146,-72.5</points>
<connection>
<GID>442</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>143.5,-59,146,-59</points>
<connection>
<GID>480</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>143.5,-46,146,-46</points>
<connection>
<GID>479</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>143.5,-85.5,146,-85.5</points>
<connection>
<GID>443</GID>
<name>IN_5</name></connection>
<intersection>143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-86.5,143,-47</points>
<intersection>-86.5 6</intersection>
<intersection>-73.5 3</intersection>
<intersection>-68.5 2</intersection>
<intersection>-60 4</intersection>
<intersection>-47 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-68.5,143,-68.5</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>143,-73.5,146,-73.5</points>
<connection>
<GID>442</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>143,-60,146,-60</points>
<connection>
<GID>480</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>143,-47,146,-47</points>
<connection>
<GID>479</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>143,-86.5,146,-86.5</points>
<connection>
<GID>443</GID>
<name>IN_4</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-87.5,142.5,-48</points>
<intersection>-87.5 5</intersection>
<intersection>-74.5 2</intersection>
<intersection>-61 3</intersection>
<intersection>-48 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>138,-74.5,146,-74.5</points>
<connection>
<GID>472</GID>
<name>OUT_3</name></connection>
<connection>
<GID>442</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>142.5,-61,146,-61</points>
<connection>
<GID>480</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142.5,-48,146,-48</points>
<connection>
<GID>479</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>142.5,-87.5,146,-87.5</points>
<connection>
<GID>443</GID>
<name>IN_3</name></connection>
<intersection>142.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-88.5,142,-49</points>
<intersection>-88.5 5</intersection>
<intersection>-76.5 2</intersection>
<intersection>-75.5 4</intersection>
<intersection>-62 3</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-49,146,-49</points>
<connection>
<GID>479</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-76.5,142,-76.5</points>
<connection>
<GID>472</GID>
<name>OUT_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>142,-62,146,-62</points>
<connection>
<GID>480</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142,-75.5,146,-75.5</points>
<connection>
<GID>442</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>142,-88.5,146,-88.5</points>
<connection>
<GID>443</GID>
<name>IN_2</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-89.5,141.5,-50</points>
<intersection>-89.5 5</intersection>
<intersection>-78.5 2</intersection>
<intersection>-76.5 4</intersection>
<intersection>-63 3</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-50,146,-50</points>
<connection>
<GID>479</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-78.5,141.5,-78.5</points>
<connection>
<GID>472</GID>
<name>OUT_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141.5,-63,146,-63</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141.5,-76.5,146,-76.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>141.5,-89.5,146,-89.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-90.5,141,-51</points>
<intersection>-90.5 5</intersection>
<intersection>-80.5 2</intersection>
<intersection>-77.5 4</intersection>
<intersection>-64 3</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-51,146,-51</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-80.5,141,-80.5</points>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>141,-64,146,-64</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>141,-77.5,146,-77.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>141,-90.5,146,-90.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-42,148,-34</points>
<intersection>-42 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-34,148,-34</points>
<connection>
<GID>474</GID>
<name>OUT_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-42,149,-42</points>
<connection>
<GID>479</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-55,148,-33</points>
<intersection>-55 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-33,148,-33</points>
<connection>
<GID>474</GID>
<name>OUT_1</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-55,149,-55</points>
<connection>
<GID>480</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-68.5,148,-32</points>
<intersection>-68.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-32,148,-32</points>
<connection>
<GID>474</GID>
<name>OUT_2</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-68.5,149,-68.5</points>
<connection>
<GID>442</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-81.5,148,-31</points>
<intersection>-81.5 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-31,148,-31</points>
<connection>
<GID>474</GID>
<name>OUT_3</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-81.5,149,-81.5</points>
<connection>
<GID>443</GID>
<name>load</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-32,132,-32</points>
<connection>
<GID>475</GID>
<name>OUT_0</name></connection>
<intersection>132 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132,-32,132,-31</points>
<connection>
<GID>474</GID>
<name>ENABLE</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-48,136.5,-37</points>
<intersection>-48 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-37,136.5,-37</points>
<intersection>131.5 3</intersection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-48,136.5,-48</points>
<connection>
<GID>477</GID>
<name>OUT_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-37,131.5,-34</points>
<intersection>-37 1</intersection>
<intersection>-34 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>131.5,-34,132,-34</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>131.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-46,137,-36.5</points>
<intersection>-46 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-36.5,137,-36.5</points>
<intersection>132 3</intersection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-46,137,-46</points>
<connection>
<GID>477</GID>
<name>OUT_1</name></connection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132,-36.5,132,-33</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire></page 4>
<page 5>
<PageViewport>-167.143,-28.8258,155.936,-199.451</PageViewport>
<gate>
<ID>582</ID>
<type>AA_LABEL</type>
<position>50.5,-56.5</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>583</ID>
<type>AA_INVERTER</type>
<position>-1.5,-21.5</position>
<input>
<ID>IN_0</ID>751 </input>
<output>
<ID>OUT_0</ID>752 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_TOGGLE</type>
<position>23,3</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_LABEL</type>
<position>0.5,-29</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>AA_LABEL</type>
<position>0.5,-30.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>587</ID>
<type>AE_REGISTER8</type>
<position>27.5,-13</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>690 </input>
<input>
<ID>IN_2</ID>691 </input>
<input>
<ID>IN_3</ID>692 </input>
<input>
<ID>IN_4</ID>693 </input>
<input>
<ID>IN_5</ID>694 </input>
<input>
<ID>IN_6</ID>695 </input>
<input>
<ID>IN_7</ID>696 </input>
<output>
<ID>OUT_0</ID>704 </output>
<output>
<ID>OUT_1</ID>703 </output>
<output>
<ID>OUT_2</ID>702 </output>
<output>
<ID>OUT_3</ID>701 </output>
<output>
<ID>OUT_4</ID>700 </output>
<output>
<ID>OUT_5</ID>699 </output>
<output>
<ID>OUT_6</ID>698 </output>
<output>
<ID>OUT_7</ID>697 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>750 </input>
<input>
<ID>count_enable</ID>712 </input>
<input>
<ID>count_up</ID>712 </input>
<input>
<ID>load</ID>752 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-72.5</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>939 </output>
<output>
<ID>OUT_1</ID>938 </output>
<output>
<ID>OUT_2</ID>937 </output>
<output>
<ID>OUT_3</ID>936 </output>
<output>
<ID>OUT_4</ID>935 </output>
<output>
<ID>OUT_5</ID>934 </output>
<output>
<ID>OUT_6</ID>933 </output>
<output>
<ID>OUT_7</ID>932 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>993 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 169</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_REGISTER8</type>
<position>44.5,-13</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>703 </input>
<input>
<ID>IN_2</ID>702 </input>
<input>
<ID>IN_3</ID>701 </input>
<input>
<ID>IN_4</ID>700 </input>
<input>
<ID>IN_5</ID>699 </input>
<input>
<ID>IN_6</ID>698 </input>
<input>
<ID>IN_7</ID>697 </input>
<output>
<ID>OUT_0</ID>715 </output>
<output>
<ID>OUT_1</ID>714 </output>
<output>
<ID>OUT_2</ID>710 </output>
<output>
<ID>OUT_3</ID>709 </output>
<output>
<ID>OUT_4</ID>708 </output>
<output>
<ID>OUT_5</ID>707 </output>
<output>
<ID>OUT_6</ID>706 </output>
<output>
<ID>OUT_7</ID>705 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>711 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-85.5</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>947 </output>
<output>
<ID>OUT_1</ID>946 </output>
<output>
<ID>OUT_2</ID>945 </output>
<output>
<ID>OUT_3</ID>944 </output>
<output>
<ID>OUT_4</ID>943 </output>
<output>
<ID>OUT_5</ID>942 </output>
<output>
<ID>OUT_6</ID>941 </output>
<output>
<ID>OUT_7</ID>940 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>994 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 147</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_REGISTER8</type>
<position>82.5,-51.5</position>
<input>
<ID>IN_0</ID>739 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>741 </input>
<input>
<ID>IN_3</ID>742 </input>
<input>
<ID>IN_4</ID>743 </input>
<input>
<ID>IN_5</ID>738 </input>
<input>
<ID>IN_6</ID>745 </input>
<input>
<ID>IN_7</ID>744 </input>
<output>
<ID>OUT_0</ID>723 </output>
<output>
<ID>OUT_1</ID>722 </output>
<output>
<ID>OUT_2</ID>721 </output>
<output>
<ID>OUT_3</ID>720 </output>
<output>
<ID>OUT_4</ID>719 </output>
<output>
<ID>OUT_5</ID>718 </output>
<output>
<ID>OUT_6</ID>717 </output>
<output>
<ID>OUT_7</ID>716 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>713 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>590</ID>
<type>AE_RAM_8x8</type>
<position>59.5,-12.5</position>
<input>
<ID>ADDRESS_0</ID>715 </input>
<input>
<ID>ADDRESS_1</ID>714 </input>
<input>
<ID>ADDRESS_2</ID>710 </input>
<input>
<ID>ADDRESS_3</ID>709 </input>
<input>
<ID>ADDRESS_4</ID>708 </input>
<input>
<ID>ADDRESS_5</ID>707 </input>
<input>
<ID>ADDRESS_6</ID>706 </input>
<input>
<ID>ADDRESS_7</ID>705 </input>
<input>
<ID>DATA_IN_0</ID>746 </input>
<input>
<ID>DATA_IN_1</ID>731 </input>
<input>
<ID>DATA_IN_2</ID>732 </input>
<input>
<ID>DATA_IN_3</ID>733 </input>
<input>
<ID>DATA_IN_4</ID>734 </input>
<input>
<ID>DATA_IN_5</ID>735 </input>
<input>
<ID>DATA_IN_6</ID>736 </input>
<input>
<ID>DATA_IN_7</ID>737 </input>
<output>
<ID>DATA_OUT_0</ID>746 </output>
<output>
<ID>DATA_OUT_1</ID>731 </output>
<output>
<ID>DATA_OUT_2</ID>732 </output>
<output>
<ID>DATA_OUT_3</ID>733 </output>
<output>
<ID>DATA_OUT_4</ID>734 </output>
<output>
<ID>DATA_OUT_5</ID>735 </output>
<output>
<ID>DATA_OUT_6</ID>736 </output>
<output>
<ID>DATA_OUT_7</ID>737 </output>
<input>
<ID>ENABLE_0</ID>730 </input>
<input>
<ID>write_enable</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>591</ID>
<type>AE_REGISTER8</type>
<position>100,-51.5</position>
<input>
<ID>IN_0</ID>723 </input>
<input>
<ID>IN_1</ID>722 </input>
<input>
<ID>IN_2</ID>721 </input>
<input>
<ID>IN_3</ID>720 </input>
<input>
<ID>IN_4</ID>719 </input>
<input>
<ID>IN_5</ID>718 </input>
<input>
<ID>IN_6</ID>717 </input>
<input>
<ID>IN_7</ID>716 </input>
<output>
<ID>OUT_0</ID>725 </output>
<output>
<ID>OUT_1</ID>726 </output>
<input>
<ID>clear</ID>728 </input>
<input>
<ID>clock</ID>727 </input>
<input>
<ID>load</ID>724 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>592</ID>
<type>DD_KEYPAD_HEX</type>
<position>8,-19</position>
<output>
<ID>OUT_0</ID>689 </output>
<output>
<ID>OUT_1</ID>690 </output>
<output>
<ID>OUT_2</ID>691 </output>
<output>
<ID>OUT_3</ID>692 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>593</ID>
<type>DD_KEYPAD_HEX</type>
<position>8,-7</position>
<output>
<ID>OUT_0</ID>693 </output>
<output>
<ID>OUT_1</ID>694 </output>
<output>
<ID>OUT_2</ID>695 </output>
<output>
<ID>OUT_3</ID>696 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>594</ID>
<type>BB_CLOCK</type>
<position>-3.5,-44.5</position>
<output>
<ID>CLK</ID>748 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>595</ID>
<type>AA_TOGGLE</type>
<position>25.5,6</position>
<output>
<ID>OUT_0</ID>712 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_LABEL</type>
<position>13,4</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>597</ID>
<type>AA_LABEL</type>
<position>13,6.5</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>598</ID>
<type>AA_TOGGLE</type>
<position>38.5,3.5</position>
<output>
<ID>OUT_0</ID>711 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_TOGGLE</type>
<position>26.5,-41.5</position>
<output>
<ID>OUT_0</ID>728 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_LABEL</type>
<position>21,-38.5</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>601</ID>
<type>AA_TOGGLE</type>
<position>79.5,-59.5</position>
<output>
<ID>OUT_0</ID>713 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>602</ID>
<type>AA_LABEL</type>
<position>22.5,-5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>603</ID>
<type>AA_LABEL</type>
<position>39,-5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>604</ID>
<type>AA_LABEL</type>
<position>59.5,-4</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>605</ID>
<type>AA_LABEL</type>
<position>86.5,-59</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>606</ID>
<type>AA_TOGGLE</type>
<position>96.5,-59.5</position>
<output>
<ID>OUT_0</ID>724 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>607</ID>
<type>BE_ROM_8x8</type>
<position>112.5,-51</position>
<input>
<ID>ADDRESS_0</ID>725 </input>
<input>
<ID>ADDRESS_1</ID>726 </input>
<input>
<ID>ENABLE_0</ID>747 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_TOGGLE</type>
<position>69.5,-10</position>
<output>
<ID>OUT_0</ID>729 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_TOGGLE</type>
<position>69.5,-13</position>
<output>
<ID>OUT_0</ID>730 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_LABEL</type>
<position>76,-9.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>611</ID>
<type>AA_LABEL</type>
<position>76.5,-12.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>612</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>73,-51</position>
<input>
<ID>ENABLE_0</ID>730 </input>
<input>
<ID>IN_0</ID>746 </input>
<input>
<ID>IN_1</ID>731 </input>
<input>
<ID>IN_2</ID>732 </input>
<input>
<ID>IN_3</ID>733 </input>
<input>
<ID>IN_4</ID>734 </input>
<input>
<ID>IN_5</ID>735 </input>
<input>
<ID>IN_6</ID>736 </input>
<input>
<ID>IN_7</ID>737 </input>
<output>
<ID>OUT_0</ID>739 </output>
<output>
<ID>OUT_1</ID>740 </output>
<output>
<ID>OUT_2</ID>741 </output>
<output>
<ID>OUT_3</ID>742 </output>
<output>
<ID>OUT_4</ID>743 </output>
<output>
<ID>OUT_5</ID>738 </output>
<output>
<ID>OUT_6</ID>745 </output>
<output>
<ID>OUT_7</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>613</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>51,-51</position>
<input>
<ID>ENABLE_0</ID>729 </input>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>962 </input>
<input>
<ID>IN_2</ID>961 </input>
<input>
<ID>IN_3</ID>960 </input>
<input>
<ID>IN_4</ID>959 </input>
<input>
<ID>IN_5</ID>958 </input>
<input>
<ID>IN_6</ID>957 </input>
<input>
<ID>IN_7</ID>956 </input>
<output>
<ID>OUT_0</ID>746 </output>
<output>
<ID>OUT_1</ID>731 </output>
<output>
<ID>OUT_2</ID>732 </output>
<output>
<ID>OUT_3</ID>733 </output>
<output>
<ID>OUT_4</ID>734 </output>
<output>
<ID>OUT_5</ID>735 </output>
<output>
<ID>OUT_6</ID>736 </output>
<output>
<ID>OUT_7</ID>737 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>614</ID>
<type>AA_LABEL</type>
<position>101.5,-58.5</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>615</ID>
<type>AA_TOGGLE</type>
<position>121.5,-30.5</position>
<output>
<ID>OUT_0</ID>747 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_LABEL</type>
<position>123,-27.5</position>
<gparam>LABEL_TEXT Output Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>22.5,-26</position>
<input>
<ID>IN_0</ID>727 </input>
<input>
<ID>IN_1</ID>751 </input>
<output>
<ID>OUT</ID>750 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_AND2</type>
<position>8,-43.5</position>
<input>
<ID>IN_0</ID>749 </input>
<input>
<ID>IN_1</ID>748 </input>
<output>
<ID>OUT</ID>727 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_TOGGLE</type>
<position>2.5,-40.5</position>
<output>
<ID>OUT_0</ID>749 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>620</ID>
<type>AA_TOGGLE</type>
<position>-6.5,-27</position>
<output>
<ID>OUT_0</ID>751 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>621</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>46.5,-85.5</position>
<input>
<ID>ENABLE_0</ID>772 </input>
<input>
<ID>IN_0</ID>1004 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1010 </input>
<input>
<ID>IN_11</ID>1017 </input>
<input>
<ID>IN_12</ID>1012 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1013 </input>
<input>
<ID>IN_15</ID>1019 </input>
<input>
<ID>IN_2</ID>1006 </input>
<input>
<ID>IN_3</ID>1007 </input>
<input>
<ID>IN_4</ID>1008 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1009 </input>
<input>
<ID>IN_7</ID>1015 </input>
<input>
<ID>IN_8</ID>1010 </input>
<input>
<ID>IN_9</ID>1016 </input>
<output>
<ID>OUT_0</ID>790 </output>
<output>
<ID>OUT_1</ID>791 </output>
<output>
<ID>OUT_10</ID>800 </output>
<output>
<ID>OUT_11</ID>801 </output>
<output>
<ID>OUT_12</ID>802 </output>
<output>
<ID>OUT_13</ID>803 </output>
<output>
<ID>OUT_14</ID>804 </output>
<output>
<ID>OUT_15</ID>805 </output>
<output>
<ID>OUT_2</ID>792 </output>
<output>
<ID>OUT_3</ID>793 </output>
<output>
<ID>OUT_4</ID>794 </output>
<output>
<ID>OUT_5</ID>795 </output>
<output>
<ID>OUT_6</ID>796 </output>
<output>
<ID>OUT_7</ID>797 </output>
<output>
<ID>OUT_8</ID>798 </output>
<output>
<ID>OUT_9</ID>799 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>622</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>46.5,-108.5</position>
<input>
<ID>ENABLE_0</ID>771 </input>
<input>
<ID>IN_0</ID>1004 </input>
<input>
<ID>IN_1</ID>1005 </input>
<input>
<ID>IN_10</ID>1011 </input>
<input>
<ID>IN_11</ID>1017 </input>
<input>
<ID>IN_12</ID>1012 </input>
<input>
<ID>IN_13</ID>1018 </input>
<input>
<ID>IN_14</ID>1013 </input>
<input>
<ID>IN_15</ID>1019 </input>
<input>
<ID>IN_2</ID>1006 </input>
<input>
<ID>IN_3</ID>1007 </input>
<input>
<ID>IN_4</ID>1008 </input>
<input>
<ID>IN_5</ID>1014 </input>
<input>
<ID>IN_6</ID>1009 </input>
<input>
<ID>IN_7</ID>1015 </input>
<input>
<ID>IN_8</ID>1010 </input>
<input>
<ID>IN_9</ID>1016 </input>
<output>
<ID>OUT_0</ID>774 </output>
<output>
<ID>OUT_1</ID>782 </output>
<output>
<ID>OUT_10</ID>779 </output>
<output>
<ID>OUT_11</ID>787 </output>
<output>
<ID>OUT_12</ID>780 </output>
<output>
<ID>OUT_13</ID>788 </output>
<output>
<ID>OUT_14</ID>781 </output>
<output>
<ID>OUT_15</ID>789 </output>
<output>
<ID>OUT_2</ID>775 </output>
<output>
<ID>OUT_3</ID>783 </output>
<output>
<ID>OUT_4</ID>776 </output>
<output>
<ID>OUT_5</ID>784 </output>
<output>
<ID>OUT_6</ID>777 </output>
<output>
<ID>OUT_7</ID>785 </output>
<output>
<ID>OUT_8</ID>778 </output>
<output>
<ID>OUT_9</ID>786 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_LABEL</type>
<position>24,-72.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>626</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-99</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>955 </output>
<output>
<ID>OUT_1</ID>954 </output>
<output>
<ID>OUT_2</ID>953 </output>
<output>
<ID>OUT_3</ID>952 </output>
<output>
<ID>OUT_4</ID>951 </output>
<output>
<ID>OUT_5</ID>950 </output>
<output>
<ID>OUT_6</ID>949 </output>
<output>
<ID>OUT_7</ID>948 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>995 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_REGISTER8</type>
<position>-75.5,-112</position>
<input>
<ID>IN_0</ID>992 </input>
<input>
<ID>IN_1</ID>991 </input>
<input>
<ID>IN_2</ID>990 </input>
<input>
<ID>IN_3</ID>989 </input>
<input>
<ID>IN_4</ID>988 </input>
<input>
<ID>IN_5</ID>987 </input>
<input>
<ID>IN_6</ID>986 </input>
<input>
<ID>IN_7</ID>985 </input>
<output>
<ID>OUT_0</ID>971 </output>
<output>
<ID>OUT_1</ID>962 </output>
<output>
<ID>OUT_2</ID>961 </output>
<output>
<ID>OUT_3</ID>960 </output>
<output>
<ID>OUT_4</ID>959 </output>
<output>
<ID>OUT_5</ID>958 </output>
<output>
<ID>OUT_6</ID>957 </output>
<output>
<ID>OUT_7</ID>956 </output>
<input>
<ID>clock</ID>972 </input>
<input>
<ID>load</ID>996 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_MUX_4x1</type>
<position>-50,-61.5</position>
<input>
<ID>IN_0</ID>956 </input>
<input>
<ID>IN_1</ID>948 </input>
<input>
<ID>IN_2</ID>940 </input>
<input>
<ID>IN_3</ID>932 </input>
<output>
<ID>OUT</ID>963 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>629</ID>
<type>AE_MUX_4x1</type>
<position>-50,-72.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>949 </input>
<input>
<ID>IN_2</ID>941 </input>
<input>
<ID>IN_3</ID>933 </input>
<output>
<ID>OUT</ID>964 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_MUX_4x1</type>
<position>-50,-83.5</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>950 </input>
<input>
<ID>IN_2</ID>942 </input>
<input>
<ID>IN_3</ID>934 </input>
<output>
<ID>OUT</ID>965 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>631</ID>
<type>AE_MUX_4x1</type>
<position>-50,-93</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>951 </input>
<input>
<ID>IN_2</ID>943 </input>
<input>
<ID>IN_3</ID>935 </input>
<output>
<ID>OUT</ID>966 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>632</ID>
<type>AE_MUX_4x1</type>
<position>-50,-104</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>952 </input>
<input>
<ID>IN_2</ID>944 </input>
<input>
<ID>IN_3</ID>936 </input>
<output>
<ID>OUT</ID>967 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>633</ID>
<type>AE_MUX_4x1</type>
<position>-50,-115</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>953 </input>
<input>
<ID>IN_2</ID>945 </input>
<input>
<ID>IN_3</ID>937 </input>
<output>
<ID>OUT</ID>968 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>634</ID>
<type>AE_MUX_4x1</type>
<position>-50,-125.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>954 </input>
<input>
<ID>IN_2</ID>946 </input>
<input>
<ID>IN_3</ID>938 </input>
<output>
<ID>OUT</ID>969 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>635</ID>
<type>AE_MUX_4x1</type>
<position>-50,-136.5</position>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>955 </input>
<input>
<ID>IN_2</ID>947 </input>
<input>
<ID>IN_3</ID>939 </input>
<output>
<ID>OUT</ID>970 </output>
<input>
<ID>SEL_0</ID>973 </input>
<input>
<ID>SEL_1</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>636</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-11.5,-94.5</position>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>969 </input>
<input>
<ID>IN_2</ID>968 </input>
<input>
<ID>IN_3</ID>967 </input>
<input>
<ID>IN_4</ID>966 </input>
<input>
<ID>IN_5</ID>965 </input>
<input>
<ID>IN_6</ID>964 </input>
<input>
<ID>IN_7</ID>963 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 147</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>637</ID>
<type>DD_KEYPAD_HEX</type>
<position>-108.5,-76.5</position>
<output>
<ID>OUT_0</ID>973 </output>
<output>
<ID>OUT_1</ID>974 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>638</ID>
<type>BB_CLOCK</type>
<position>-87,-120.5</position>
<output>
<ID>CLK</ID>972 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_LABEL</type>
<position>-75,-105</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>640</ID>
<type>AA_LABEL</type>
<position>-75,-91.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>641</ID>
<type>AA_LABEL</type>
<position>-75,-78.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>642</ID>
<type>AA_LABEL</type>
<position>-75,-65</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>643</ID>
<type>AA_LABEL</type>
<position>-110,-69.5</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>644</ID>
<type>DD_KEYPAD_HEX</type>
<position>-108.5,-90.5</position>
<output>
<ID>OUT_0</ID>983 </output>
<output>
<ID>OUT_1</ID>984 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-61.5</position>
<input>
<ID>IN_0</ID>932 </input>
<input>
<ID>IN_1</ID>948 </input>
<input>
<ID>IN_2</ID>940 </input>
<input>
<ID>IN_3</ID>932 </input>
<output>
<ID>OUT</ID>975 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-72.5</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>949 </input>
<input>
<ID>IN_2</ID>941 </input>
<input>
<ID>IN_3</ID>933 </input>
<output>
<ID>OUT</ID>976 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-83.5</position>
<input>
<ID>IN_0</ID>958 </input>
<input>
<ID>IN_1</ID>950 </input>
<input>
<ID>IN_2</ID>942 </input>
<input>
<ID>IN_3</ID>934 </input>
<output>
<ID>OUT</ID>977 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>648</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-93</position>
<input>
<ID>IN_0</ID>959 </input>
<input>
<ID>IN_1</ID>951 </input>
<input>
<ID>IN_2</ID>943 </input>
<input>
<ID>IN_3</ID>935 </input>
<output>
<ID>OUT</ID>978 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-104</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>952 </input>
<input>
<ID>IN_2</ID>944 </input>
<input>
<ID>IN_3</ID>936 </input>
<output>
<ID>OUT</ID>979 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-115</position>
<input>
<ID>IN_0</ID>961 </input>
<input>
<ID>IN_1</ID>953 </input>
<input>
<ID>IN_2</ID>945 </input>
<input>
<ID>IN_3</ID>937 </input>
<output>
<ID>OUT</ID>980 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>651</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-125.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>954 </input>
<input>
<ID>IN_2</ID>946 </input>
<input>
<ID>IN_3</ID>938 </input>
<output>
<ID>OUT</ID>981 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>652</ID>
<type>AE_MUX_4x1</type>
<position>-37.5,-136.5</position>
<input>
<ID>IN_0</ID>971 </input>
<input>
<ID>IN_1</ID>955 </input>
<input>
<ID>IN_2</ID>947 </input>
<input>
<ID>IN_3</ID>939 </input>
<output>
<ID>OUT</ID>982 </output>
<input>
<ID>SEL_0</ID>983 </input>
<input>
<ID>SEL_1</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>653</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-9.5,-105</position>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>980 </input>
<input>
<ID>IN_3</ID>979 </input>
<input>
<ID>IN_4</ID>978 </input>
<input>
<ID>IN_5</ID>977 </input>
<input>
<ID>IN_6</ID>976 </input>
<input>
<ID>IN_7</ID>975 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 169</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>654</ID>
<type>AA_LABEL</type>
<position>-110,-83.5</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>655</ID>
<type>DD_KEYPAD_HEX</type>
<position>-92.5,-90</position>
<output>
<ID>OUT_0</ID>988 </output>
<output>
<ID>OUT_1</ID>987 </output>
<output>
<ID>OUT_2</ID>986 </output>
<output>
<ID>OUT_3</ID>985 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 9</lparam></gate>
<gate>
<ID>656</ID>
<type>DD_KEYPAD_HEX</type>
<position>-92.5,-102</position>
<output>
<ID>OUT_0</ID>992 </output>
<output>
<ID>OUT_1</ID>991 </output>
<output>
<ID>OUT_2</ID>990 </output>
<output>
<ID>OUT_3</ID>989 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_LABEL</type>
<position>-92.5,-83</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>658</ID>
<type>BA_DECODER_2x4</type>
<position>-90.5,-57</position>
<input>
<ID>ENABLE</ID>997 </input>
<input>
<ID>IN_0</ID>998 </input>
<input>
<ID>IN_1</ID>999 </input>
<output>
<ID>OUT_0</ID>993 </output>
<output>
<ID>OUT_1</ID>994 </output>
<output>
<ID>OUT_2</ID>995 </output>
<output>
<ID>OUT_3</ID>996 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_TOGGLE</type>
<position>-96.5,-56.5</position>
<output>
<ID>OUT_0</ID>997 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_LABEL</type>
<position>-99,-55</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>661</ID>
<type>DD_KEYPAD_HEX</type>
<position>-95.5,-69.5</position>
<output>
<ID>OUT_0</ID>998 </output>
<output>
<ID>OUT_1</ID>999 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_LABEL</type>
<position>-95,-62.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>668</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>6.5,-83.5</position>
<input>
<ID>ENABLE_0</ID>1000 </input>
<input>
<ID>IN_0</ID>970 </input>
<input>
<ID>IN_1</ID>969 </input>
<input>
<ID>IN_2</ID>968 </input>
<input>
<ID>IN_3</ID>967 </input>
<input>
<ID>IN_4</ID>966 </input>
<input>
<ID>IN_5</ID>965 </input>
<input>
<ID>IN_6</ID>964 </input>
<input>
<ID>IN_7</ID>963 </input>
<output>
<ID>OUT_0</ID>1005 </output>
<output>
<ID>OUT_1</ID>1007 </output>
<output>
<ID>OUT_2</ID>1014 </output>
<output>
<ID>OUT_3</ID>1015 </output>
<output>
<ID>OUT_4</ID>1016 </output>
<output>
<ID>OUT_5</ID>1017 </output>
<output>
<ID>OUT_6</ID>1018 </output>
<output>
<ID>OUT_7</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>670</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>6.5,-115</position>
<input>
<ID>ENABLE_0</ID>1002 </input>
<input>
<ID>IN_0</ID>982 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>980 </input>
<input>
<ID>IN_3</ID>979 </input>
<input>
<ID>IN_4</ID>978 </input>
<input>
<ID>IN_5</ID>977 </input>
<input>
<ID>IN_6</ID>976 </input>
<input>
<ID>IN_7</ID>975 </input>
<output>
<ID>OUT_0</ID>1004 </output>
<output>
<ID>OUT_1</ID>1006 </output>
<output>
<ID>OUT_2</ID>1008 </output>
<output>
<ID>OUT_3</ID>1009 </output>
<output>
<ID>OUT_4</ID>1010 </output>
<output>
<ID>OUT_5</ID>1011 </output>
<output>
<ID>OUT_6</ID>1012 </output>
<output>
<ID>OUT_7</ID>1013 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>672</ID>
<type>EE_VDD</type>
<position>6.5,-71.5</position>
<output>
<ID>OUT_0</ID>1000 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_LABEL</type>
<position>4,-74.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>482</ID>
<type>AA_LABEL</type>
<position>-18.5,-88</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>676</ID>
<type>AA_LABEL</type>
<position>6.5,-121</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>484</ID>
<type>AA_LABEL</type>
<position>-18.5,-99</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>678</ID>
<type>EE_VDD</type>
<position>6.5,-100</position>
<output>
<ID>OUT_0</ID>1002 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>492</ID>
<type>BA_DECODER_2x4</type>
<position>38,-69</position>
<input>
<ID>ENABLE</ID>769 </input>
<input>
<ID>IN_0</ID>770 </input>
<output>
<ID>OUT_0</ID>771 </output>
<output>
<ID>OUT_1</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_TOGGLE</type>
<position>33,-67.5</position>
<output>
<ID>OUT_0</ID>769 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_TOGGLE</type>
<position>28.5,-70.5</position>
<output>
<ID>OUT_0</ID>770 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_LABEL</type>
<position>33.5,-64.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>496</ID>
<type>AA_LABEL</type>
<position>22,-70</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>497</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64,-104.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>783 </input>
<input>
<ID>IN_2</ID>784 </input>
<input>
<ID>IN_3</ID>785 </input>
<input>
<ID>IN_B_0</ID>774 </input>
<input>
<ID>IN_B_1</ID>775 </input>
<input>
<ID>IN_B_2</ID>776 </input>
<input>
<ID>IN_B_3</ID>777 </input>
<output>
<ID>OUT_0</ID>806 </output>
<output>
<ID>OUT_1</ID>807 </output>
<output>
<ID>OUT_2</ID>808 </output>
<output>
<ID>OUT_3</ID>809 </output>
<output>
<ID>carry_out</ID>773 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_FULLADDER_4BIT</type>
<position>64,-120.5</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>787 </input>
<input>
<ID>IN_2</ID>788 </input>
<input>
<ID>IN_3</ID>789 </input>
<input>
<ID>IN_B_0</ID>778 </input>
<input>
<ID>IN_B_1</ID>779 </input>
<input>
<ID>IN_B_2</ID>780 </input>
<input>
<ID>IN_B_3</ID>781 </input>
<output>
<ID>OUT_0</ID>810 </output>
<output>
<ID>OUT_1</ID>811 </output>
<output>
<ID>OUT_2</ID>812 </output>
<output>
<ID>OUT_3</ID>813 </output>
<input>
<ID>carry_in</ID>773 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_LABEL</type>
<position>71.5,-97</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>500</ID>
<type>AA_LABEL</type>
<position>72,-125.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>501</ID>
<type>AA_LABEL</type>
<position>57.5,-98</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>502</ID>
<type>AA_LABEL</type>
<position>58,-104.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>503</ID>
<type>AA_LABEL</type>
<position>57.5,-114</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>504</ID>
<type>AA_LABEL</type>
<position>58.5,-121</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>AA_AND2</type>
<position>59.5,-94</position>
<input>
<ID>IN_0</ID>791 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_AND2</type>
<position>64.5,-90.5</position>
<input>
<ID>IN_0</ID>793 </input>
<input>
<ID>IN_1</ID>792 </input>
<output>
<ID>OUT</ID>815 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_AND2</type>
<position>59.5,-87</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>794 </input>
<output>
<ID>OUT</ID>816 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_AND2</type>
<position>64.5,-83.5</position>
<input>
<ID>IN_0</ID>797 </input>
<input>
<ID>IN_1</ID>796 </input>
<output>
<ID>OUT</ID>817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>59.5,-80</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>798 </input>
<output>
<ID>OUT</ID>818 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_AND2</type>
<position>64.5,-76.5</position>
<input>
<ID>IN_0</ID>801 </input>
<input>
<ID>IN_1</ID>800 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_AND2</type>
<position>59.5,-73</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>802 </input>
<output>
<ID>OUT</ID>820 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>64.5,-69.5</position>
<input>
<ID>IN_0</ID>805 </input>
<input>
<ID>IN_1</ID>804 </input>
<output>
<ID>OUT</ID>821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-81</position>
<input>
<ID>IN_0</ID>813 </input>
<input>
<ID>IN_1</ID>821 </input>
<output>
<ID>OUT</ID>829 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-86</position>
<input>
<ID>IN_0</ID>812 </input>
<input>
<ID>IN_1</ID>820 </input>
<output>
<ID>OUT</ID>828 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-91</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>819 </input>
<output>
<ID>OUT</ID>827 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-96</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>818 </input>
<output>
<ID>OUT</ID>826 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>517</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-101</position>
<input>
<ID>IN_0</ID>809 </input>
<input>
<ID>IN_1</ID>817 </input>
<output>
<ID>OUT</ID>825 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-106</position>
<input>
<ID>IN_0</ID>808 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>824 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-111</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>815 </input>
<output>
<ID>OUT</ID>823 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AA_MUX_2x1</type>
<position>89.5,-116</position>
<input>
<ID>IN_0</ID>806 </input>
<input>
<ID>IN_1</ID>814 </input>
<output>
<ID>OUT</ID>822 </output>
<input>
<ID>SEL_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>521</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>112,-98</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>823 </input>
<input>
<ID>IN_2</ID>824 </input>
<input>
<ID>IN_3</ID>825 </input>
<input>
<ID>IN_4</ID>826 </input>
<input>
<ID>IN_5</ID>827 </input>
<input>
<ID>IN_6</ID>828 </input>
<input>
<ID>IN_7</ID>829 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 60</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_LABEL</type>
<position>89.5,-119.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>523</ID>
<type>AA_LABEL</type>
<position>90.5,-77</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>524</ID>
<type>GA_LED</type>
<position>103.5,-108</position>
<input>
<ID>N_in2</ID>829 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>525</ID>
<type>GA_LED</type>
<position>106,-108</position>
<input>
<ID>N_in2</ID>828 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>526</ID>
<type>GA_LED</type>
<position>108.5,-108</position>
<input>
<ID>N_in2</ID>827 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>527</ID>
<type>GA_LED</type>
<position>111,-108</position>
<input>
<ID>N_in2</ID>826 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>528</ID>
<type>GA_LED</type>
<position>113.5,-108</position>
<input>
<ID>N_in2</ID>825 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>529</ID>
<type>GA_LED</type>
<position>116,-108</position>
<input>
<ID>N_in2</ID>824 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>530</ID>
<type>GA_LED</type>
<position>118.5,-108</position>
<input>
<ID>N_in2</ID>823 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>531</ID>
<type>GA_LED</type>
<position>121,-108</position>
<input>
<ID>N_in2</ID>822 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>532</ID>
<type>AA_LABEL</type>
<position>121,-110</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>533</ID>
<type>AA_LABEL</type>
<position>118.5,-110</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>534</ID>
<type>AA_LABEL</type>
<position>116,-110</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>535</ID>
<type>AA_LABEL</type>
<position>113.5,-110</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>536</ID>
<type>AA_LABEL</type>
<position>111,-110</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>537</ID>
<type>AA_LABEL</type>
<position>108.5,-110</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>AA_LABEL</type>
<position>106,-110</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>539</ID>
<type>AA_LABEL</type>
<position>103.5,-110</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-115.5,53.5,-108</points>
<intersection>-115.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-115.5,60,-115.5</points>
<connection>
<GID>498</GID>
<name>IN_B_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-108,53.5,-108</points>
<connection>
<GID>622</GID>
<name>OUT_8</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-116.5,53,-106</points>
<intersection>-116.5 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-116.5,60,-116.5</points>
<connection>
<GID>498</GID>
<name>IN_B_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-106,53,-106</points>
<connection>
<GID>622</GID>
<name>OUT_10</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-117.5,52.5,-104</points>
<intersection>-117.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-117.5,60,-117.5</points>
<connection>
<GID>498</GID>
<name>IN_B_2</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-104,52.5,-104</points>
<connection>
<GID>622</GID>
<name>OUT_12</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-118.5,52,-102</points>
<intersection>-118.5 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-118.5,60,-118.5</points>
<connection>
<GID>498</GID>
<name>IN_B_3</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-102,52,-102</points>
<connection>
<GID>622</GID>
<name>OUT_14</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-115,54,-106.5</points>
<intersection>-115 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-106.5,60,-106.5</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-115,54,-115</points>
<connection>
<GID>622</GID>
<name>OUT_1</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-113,54,-107.5</points>
<intersection>-113 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-107.5,60,-107.5</points>
<connection>
<GID>497</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-113,54,-113</points>
<connection>
<GID>622</GID>
<name>OUT_3</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-111,54,-108.5</points>
<intersection>-111 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-108.5,60,-108.5</points>
<connection>
<GID>497</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-111,54,-111</points>
<connection>
<GID>622</GID>
<name>OUT_5</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-109.5,54,-109</points>
<intersection>-109.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-109.5,60,-109.5</points>
<connection>
<GID>497</GID>
<name>IN_3</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-109,54,-109</points>
<connection>
<GID>622</GID>
<name>OUT_7</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-122.5,56,-107</points>
<intersection>-122.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-122.5,60,-122.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-107,56,-107</points>
<connection>
<GID>622</GID>
<name>OUT_9</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-123.5,55.5,-105</points>
<intersection>-123.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-123.5,60,-123.5</points>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-105,55.5,-105</points>
<connection>
<GID>622</GID>
<name>OUT_11</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-124.5,55,-103</points>
<intersection>-124.5 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-124.5,60,-124.5</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-103,55,-103</points>
<connection>
<GID>622</GID>
<name>OUT_13</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-125.5,54.5,-101</points>
<intersection>-125.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-125.5,60,-125.5</points>
<connection>
<GID>498</GID>
<name>IN_3</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-101,54.5,-101</points>
<connection>
<GID>622</GID>
<name>OUT_15</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-95,49.5,-93</points>
<intersection>-95 1</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-95,56.5,-95</points>
<connection>
<GID>505</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-93,49.5,-93</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-93,56.5,-93</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-93,48.5,-92</points>
<connection>
<GID>621</GID>
<name>OUT_1</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-91.5,52,-91</points>
<intersection>-91.5 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-91.5,61.5,-91.5</points>
<connection>
<GID>506</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-91,52,-91</points>
<connection>
<GID>621</GID>
<name>OUT_2</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-89.5,61.5,-89.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-90,48.5,-89.5</points>
<connection>
<GID>621</GID>
<name>OUT_3</name></connection>
<intersection>-89.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-88,56.5,-88</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-89,48.5,-88</points>
<connection>
<GID>621</GID>
<name>OUT_4</name></connection>
<intersection>-88 1</intersection></vsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-88,49.5,-86</points>
<intersection>-88 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-86,56.5,-86</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-88,49.5,-88</points>
<connection>
<GID>621</GID>
<name>OUT_5</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-87,50.5,-84.5</points>
<intersection>-87 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-84.5,61.5,-84.5</points>
<connection>
<GID>508</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-87,50.5,-87</points>
<connection>
<GID>621</GID>
<name>OUT_6</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-86,50,-82.5</points>
<intersection>-86 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-82.5,61.5,-82.5</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-86,50,-86</points>
<connection>
<GID>621</GID>
<name>OUT_7</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-85,49.5,-81</points>
<intersection>-85 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-81,56.5,-81</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-85,49.5,-85</points>
<connection>
<GID>621</GID>
<name>OUT_8</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-84,49.5,-79</points>
<intersection>-84 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-79,56.5,-79</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-84,49.5,-84</points>
<connection>
<GID>621</GID>
<name>OUT_9</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-83,50,-77.5</points>
<intersection>-83 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-77.5,61.5,-77.5</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-83,50,-83</points>
<connection>
<GID>621</GID>
<name>OUT_10</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-82,50,-75.5</points>
<intersection>-82 2</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-75.5,61.5,-75.5</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-82,50,-82</points>
<connection>
<GID>621</GID>
<name>OUT_11</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-81,49.5,-74</points>
<intersection>-81 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-74,56.5,-74</points>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-81,49.5,-81</points>
<connection>
<GID>621</GID>
<name>OUT_12</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-80,49.5,-72</points>
<intersection>-80 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-72,56.5,-72</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-80,49.5,-80</points>
<connection>
<GID>621</GID>
<name>OUT_13</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-79,49,-70.5</points>
<intersection>-79 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-70.5,61.5,-70.5</points>
<connection>
<GID>512</GID>
<name>IN_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-79,49,-79</points>
<connection>
<GID>621</GID>
<name>OUT_14</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-78,48.5,-68.5</points>
<connection>
<GID>621</GID>
<name>OUT_15</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-68.5,61.5,-68.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-117,77.5,-103</points>
<intersection>-117 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-117,87.5,-117</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-103,77.5,-103</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-112,77.5,-104</points>
<intersection>-112 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-112,87.5,-112</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-104,77.5,-104</points>
<connection>
<GID>497</GID>
<name>OUT_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-107,77.5,-105</points>
<intersection>-107 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-107,87.5,-107</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-105,77.5,-105</points>
<connection>
<GID>497</GID>
<name>OUT_2</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-106,77.5,-102</points>
<intersection>-106 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-102,87.5,-102</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-106,77.5,-106</points>
<connection>
<GID>497</GID>
<name>OUT_3</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-119,77.5,-97</points>
<intersection>-119 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-97,87.5,-97</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-119,77.5,-119</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-120,77.5,-92</points>
<intersection>-120 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-92,87.5,-92</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-120,77.5,-120</points>
<connection>
<GID>498</GID>
<name>OUT_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-121,77.5,-87</points>
<intersection>-121 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-87,87.5,-87</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-121,77.5,-121</points>
<connection>
<GID>498</GID>
<name>OUT_2</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>813</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-122,77.5,-82</points>
<intersection>-122 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-82,87.5,-82</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-122,77.5,-122</points>
<connection>
<GID>498</GID>
<name>OUT_3</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>814</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-115,75,-94</points>
<intersection>-115 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-115,87.5,-115</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-94,75,-94</points>
<connection>
<GID>505</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>815</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-110,77.5,-90.5</points>
<intersection>-110 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-90.5,77.5,-90.5</points>
<connection>
<GID>506</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-110,87.5,-110</points>
<connection>
<GID>519</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>816</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-105,75,-87</points>
<intersection>-105 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-87,75,-87</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-105,87.5,-105</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>817</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-100,77.5,-83.5</points>
<intersection>-100 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-83.5,77.5,-83.5</points>
<connection>
<GID>508</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-100,87.5,-100</points>
<connection>
<GID>517</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-95,75,-80</points>
<intersection>-95 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-80,75,-80</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-95,87.5,-95</points>
<connection>
<GID>516</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-90,77.5,-76.5</points>
<intersection>-90 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-76.5,77.5,-76.5</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-90,87.5,-90</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-85,75,-73</points>
<intersection>-85 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-73,75,-73</points>
<connection>
<GID>511</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-85,87.5,-85</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-80,77.5,-69.5</points>
<intersection>-80 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-69.5,77.5,-69.5</points>
<connection>
<GID>512</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-80,87.5,-80</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-116,99,-101</points>
<intersection>-116 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-101,107,-101</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection>
<intersection>100 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-116,99,-116</points>
<connection>
<GID>520</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>100,-106.5,100,-101</points>
<intersection>-106.5 8</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100,-106.5,121,-106.5</points>
<intersection>100 7</intersection>
<intersection>121 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>121,-107,121,-106.5</points>
<connection>
<GID>531</GID>
<name>N_in2</name></connection>
<intersection>-106.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-111,99,-100</points>
<intersection>-111 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-100,107,-100</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection>
<intersection>100.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-111,99,-111</points>
<connection>
<GID>519</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>100.5,-106,100.5,-100</points>
<intersection>-106 8</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100.5,-106,118.5,-106</points>
<intersection>100.5 7</intersection>
<intersection>118.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>118.5,-107,118.5,-106</points>
<connection>
<GID>530</GID>
<name>N_in2</name></connection>
<intersection>-106 8</intersection></vsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-106,99,-99</points>
<intersection>-106 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-99,107,-99</points>
<connection>
<GID>521</GID>
<name>IN_2</name></connection>
<intersection>99 0</intersection>
<intersection>101 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-106,99,-106</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>101,-105.5,101,-99</points>
<intersection>-105.5 8</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>101,-105.5,116,-105.5</points>
<intersection>101 7</intersection>
<intersection>116 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>116,-107,116,-105.5</points>
<connection>
<GID>529</GID>
<name>N_in2</name></connection>
<intersection>-105.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-101,99,-98</points>
<intersection>-101 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-98,107,-98</points>
<connection>
<GID>521</GID>
<name>IN_3</name></connection>
<intersection>99 0</intersection>
<intersection>101.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-101,99,-101</points>
<connection>
<GID>517</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>101.5,-105,101.5,-98</points>
<intersection>-105 9</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>101.5,-105,113.5,-105</points>
<intersection>101.5 8</intersection>
<intersection>113.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>113.5,-107,113.5,-105</points>
<connection>
<GID>528</GID>
<name>N_in2</name></connection>
<intersection>-105 9</intersection></vsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-97,99,-96</points>
<intersection>-97 1</intersection>
<intersection>-96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-97,107,-97</points>
<connection>
<GID>521</GID>
<name>IN_4</name></connection>
<intersection>99 0</intersection>
<intersection>102 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-96,99,-96</points>
<connection>
<GID>516</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>102,-104.5,102,-97</points>
<intersection>-104.5 9</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>102,-104.5,111,-104.5</points>
<intersection>102 8</intersection>
<intersection>111 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>111,-107,111,-104.5</points>
<connection>
<GID>527</GID>
<name>N_in2</name></connection>
<intersection>-104.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-96,99,-91</points>
<intersection>-96 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-96,107,-96</points>
<connection>
<GID>521</GID>
<name>IN_5</name></connection>
<intersection>99 0</intersection>
<intersection>102.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-91,99,-91</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>102.5,-104,102.5,-96</points>
<intersection>-104 8</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>102.5,-104,108.5,-104</points>
<intersection>102.5 7</intersection>
<intersection>108.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>108.5,-107,108.5,-104</points>
<connection>
<GID>526</GID>
<name>N_in2</name></connection>
<intersection>-104 8</intersection></vsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-95,99,-86</points>
<intersection>-95 1</intersection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-95,107,-95</points>
<connection>
<GID>521</GID>
<name>IN_6</name></connection>
<intersection>99 0</intersection>
<intersection>103 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-86,99,-86</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>103,-103.5,103,-95</points>
<intersection>-103.5 8</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>103,-103.5,106,-103.5</points>
<intersection>103 7</intersection>
<intersection>106 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>106,-107,106,-103.5</points>
<connection>
<GID>525</GID>
<name>N_in2</name></connection>
<intersection>-103.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-94,99,-81</points>
<intersection>-94 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-81,99,-81</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-94,107,-94</points>
<connection>
<GID>521</GID>
<name>IN_7</name></connection>
<intersection>99 0</intersection>
<intersection>103.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>103.5,-107,103.5,-94</points>
<connection>
<GID>524</GID>
<name>N_in2</name></connection>
<intersection>-94 2</intersection></vsegment></shape></wire>
<wire>
<ID>932</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-68.5,-53.5,-68.5</points>
<connection>
<GID>202</GID>
<name>OUT_7</name></connection>
<intersection>-53.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-53.5,-68.5,-53.5,-58.5</points>
<intersection>-68.5 1</intersection>
<intersection>-58.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-53.5,-58.5,-40.5,-58.5</points>
<connection>
<GID>628</GID>
<name>IN_3</name></connection>
<connection>
<GID>645</GID>
<name>IN_3</name></connection>
<intersection>-53.5 4</intersection>
<intersection>-42 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-42,-64.5,-42,-58.5</points>
<intersection>-64.5 8</intersection>
<intersection>-58.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-42,-64.5,-40.5,-64.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>-42 6</intersection></hsegment></shape></wire>
<wire>
<ID>933</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-69.5,-40.5,-69.5</points>
<connection>
<GID>202</GID>
<name>OUT_6</name></connection>
<connection>
<GID>629</GID>
<name>IN_3</name></connection>
<connection>
<GID>646</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>934</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-80.5,-54.5,-70.5</points>
<intersection>-80.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,-80.5,-40.5,-80.5</points>
<connection>
<GID>630</GID>
<name>IN_3</name></connection>
<connection>
<GID>647</GID>
<name>IN_3</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-70.5,-54.5,-70.5</points>
<connection>
<GID>202</GID>
<name>OUT_5</name></connection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>935</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-90,-55,-71.5</points>
<intersection>-90 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-90,-40.5,-90</points>
<connection>
<GID>631</GID>
<name>IN_3</name></connection>
<connection>
<GID>648</GID>
<name>IN_3</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-71.5,-55,-71.5</points>
<connection>
<GID>202</GID>
<name>OUT_4</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-101,-55.5,-72.5</points>
<intersection>-101 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-101,-40.5,-101</points>
<connection>
<GID>632</GID>
<name>IN_3</name></connection>
<connection>
<GID>649</GID>
<name>IN_3</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-72.5,-55.5,-72.5</points>
<connection>
<GID>202</GID>
<name>OUT_3</name></connection>
<intersection>-55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-112,-56,-73.5</points>
<intersection>-112 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-112,-40.5,-112</points>
<connection>
<GID>633</GID>
<name>IN_3</name></connection>
<connection>
<GID>650</GID>
<name>IN_3</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-73.5,-56,-73.5</points>
<connection>
<GID>202</GID>
<name>OUT_2</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-122.5,-56.5,-74.5</points>
<intersection>-122.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,-122.5,-40.5,-122.5</points>
<connection>
<GID>634</GID>
<name>IN_3</name></connection>
<connection>
<GID>651</GID>
<name>IN_3</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-74.5,-56.5,-74.5</points>
<connection>
<GID>202</GID>
<name>OUT_1</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>939</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-133.5,-57,-75.5</points>
<intersection>-133.5 2</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-75.5,-57,-75.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-133.5,-40.5,-133.5</points>
<connection>
<GID>635</GID>
<name>IN_3</name></connection>
<connection>
<GID>652</GID>
<name>IN_3</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-81.5,-58,-60.5</points>
<intersection>-81.5 2</intersection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-60.5,-40.5,-60.5</points>
<connection>
<GID>628</GID>
<name>IN_2</name></connection>
<connection>
<GID>645</GID>
<name>IN_2</name></connection>
<intersection>-58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-81.5,-58,-81.5</points>
<connection>
<GID>203</GID>
<name>OUT_7</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>941</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-82.5,-58.5,-71.5</points>
<intersection>-82.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-71.5,-40.5,-71.5</points>
<connection>
<GID>629</GID>
<name>IN_2</name></connection>
<connection>
<GID>646</GID>
<name>IN_2</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-82.5,-58.5,-82.5</points>
<connection>
<GID>203</GID>
<name>OUT_6</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>942</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71.5,-83.5,-53,-83.5</points>
<connection>
<GID>203</GID>
<name>OUT_5</name></connection>
<intersection>-53 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-53,-83.5,-53,-82.5</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>-83.5 1</intersection>
<intersection>-82.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-53,-82.5,-40.5,-82.5</points>
<connection>
<GID>647</GID>
<name>IN_2</name></connection>
<intersection>-53 3</intersection></hsegment></shape></wire>
<wire>
<ID>943</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-92,-59,-84.5</points>
<intersection>-92 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,-92,-40.5,-92</points>
<connection>
<GID>631</GID>
<name>IN_2</name></connection>
<connection>
<GID>648</GID>
<name>IN_2</name></connection>
<intersection>-59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-84.5,-59,-84.5</points>
<connection>
<GID>203</GID>
<name>OUT_4</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-103,-59.5,-85.5</points>
<intersection>-103 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-103,-40.5,-103</points>
<connection>
<GID>632</GID>
<name>IN_2</name></connection>
<connection>
<GID>649</GID>
<name>IN_2</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-85.5,-59.5,-85.5</points>
<connection>
<GID>203</GID>
<name>OUT_3</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>945</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-114,-60,-86.5</points>
<intersection>-114 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-114,-40.5,-114</points>
<connection>
<GID>633</GID>
<name>IN_2</name></connection>
<connection>
<GID>650</GID>
<name>IN_2</name></connection>
<intersection>-60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-86.5,-60,-86.5</points>
<connection>
<GID>203</GID>
<name>OUT_2</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>946</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-124.5,-60.5,-87.5</points>
<intersection>-124.5 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-87.5,-60.5,-87.5</points>
<connection>
<GID>203</GID>
<name>OUT_1</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-60.5,-124.5,-40.5,-124.5</points>
<connection>
<GID>634</GID>
<name>IN_2</name></connection>
<connection>
<GID>651</GID>
<name>IN_2</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>947</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-135.5,-57.5,-88.5</points>
<intersection>-135.5 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,-135.5,-40.5,-135.5</points>
<connection>
<GID>635</GID>
<name>IN_2</name></connection>
<connection>
<GID>652</GID>
<name>IN_2</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-88.5,-57.5,-88.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-95,-62,-62.5</points>
<intersection>-95 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-62.5,-40.5,-62.5</points>
<connection>
<GID>628</GID>
<name>IN_1</name></connection>
<connection>
<GID>645</GID>
<name>IN_1</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-95,-62,-95</points>
<connection>
<GID>626</GID>
<name>OUT_7</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-96,-62.5,-73.5</points>
<intersection>-96 2</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-73.5,-40.5,-73.5</points>
<connection>
<GID>629</GID>
<name>IN_1</name></connection>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-96,-62.5,-96</points>
<connection>
<GID>626</GID>
<name>OUT_6</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>950</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-97,-63,-84.5</points>
<intersection>-97 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-84.5,-40.5,-84.5</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<connection>
<GID>647</GID>
<name>IN_1</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-97,-63,-97</points>
<connection>
<GID>626</GID>
<name>OUT_5</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-98,-63.5,-94</points>
<intersection>-98 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-94,-40.5,-94</points>
<connection>
<GID>631</GID>
<name>IN_1</name></connection>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-98,-63.5,-98</points>
<connection>
<GID>626</GID>
<name>OUT_4</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>952</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,-105,-64,-99</points>
<intersection>-105 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-105,-40.5,-105</points>
<connection>
<GID>632</GID>
<name>IN_1</name></connection>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-99,-64,-99</points>
<connection>
<GID>626</GID>
<name>OUT_3</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>953</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-116,-64.5,-100</points>
<intersection>-116 1</intersection>
<intersection>-100 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-116,-40.5,-116</points>
<connection>
<GID>633</GID>
<name>IN_1</name></connection>
<connection>
<GID>650</GID>
<name>IN_1</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-100,-64.5,-100</points>
<connection>
<GID>626</GID>
<name>OUT_2</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-126.5,-65,-101</points>
<intersection>-126.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-126.5,-40.5,-126.5</points>
<connection>
<GID>634</GID>
<name>IN_1</name></connection>
<connection>
<GID>651</GID>
<name>IN_1</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-101,-65,-101</points>
<connection>
<GID>626</GID>
<name>OUT_1</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>955</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-137.5,-65.5,-102</points>
<intersection>-137.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71.5,-102,-65.5,-102</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,-137.5,-40.5,-137.5</points>
<connection>
<GID>635</GID>
<name>IN_1</name></connection>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-153,-66.5,-108</points>
<intersection>-153 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,-153,-4.5,-153</points>
<intersection>-66.5 0</intersection>
<intersection>-53 5</intersection>
<intersection>-4.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-108,-66.5,-108</points>
<connection>
<GID>627</GID>
<name>OUT_7</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-4.5,-153,-4.5,-47.5</points>
<intersection>-153 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-53,-153,-53,-64.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-4.5,-47.5,49,-47.5</points>
<connection>
<GID>613</GID>
<name>IN_7</name></connection>
<intersection>-4.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>957</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,-154.5,-67,-109</points>
<intersection>-154.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,-154.5,-3,-154.5</points>
<intersection>-67 0</intersection>
<intersection>-53 7</intersection>
<intersection>-40.5 8</intersection>
<intersection>-3 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-109,-67,-109</points>
<connection>
<GID>627</GID>
<name>OUT_6</name></connection>
<intersection>-67 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-3,-154.5,-3,-48.5</points>
<intersection>-154.5 1</intersection>
<intersection>-48.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-3,-48.5,49,-48.5</points>
<connection>
<GID>613</GID>
<name>IN_6</name></connection>
<intersection>-3 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-53,-154.5,-53,-75.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-40.5,-154.5,-40.5,-75.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>958</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-155.5,-67.5,-110</points>
<intersection>-155.5 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67.5,-155.5,-1.5,-155.5</points>
<intersection>-67.5 0</intersection>
<intersection>-53 8</intersection>
<intersection>-40.5 9</intersection>
<intersection>-1.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-110,-67.5,-110</points>
<connection>
<GID>627</GID>
<name>OUT_5</name></connection>
<intersection>-67.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-1.5,-155.5,-1.5,-49.5</points>
<intersection>-155.5 1</intersection>
<intersection>-49.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-1.5,-49.5,49,-49.5</points>
<connection>
<GID>613</GID>
<name>IN_5</name></connection>
<intersection>-1.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-53,-155.5,-53,-86.5</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>-155.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-40.5,-155.5,-40.5,-86.5</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-155.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-157.5,0,-157.5</points>
<intersection>-68 6</intersection>
<intersection>-53 13</intersection>
<intersection>-40.5 14</intersection>
<intersection>0 11</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-68,-157.5,-68,-111</points>
<intersection>-157.5 1</intersection>
<intersection>-111 15</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>0,-157.5,0,-50.5</points>
<intersection>-157.5 1</intersection>
<intersection>-50.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>0,-50.5,49,-50.5</points>
<connection>
<GID>613</GID>
<name>IN_4</name></connection>
<intersection>0 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-53,-157.5,-53,-96</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-40.5,-157.5,-40.5,-96</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-71.5,-111,-68,-111</points>
<connection>
<GID>627</GID>
<name>OUT_4</name></connection>
<intersection>-68 6</intersection></hsegment></shape></wire>
<wire>
<ID>960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-159,-68.5,-112</points>
<intersection>-159 1</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,-159,1,-159</points>
<intersection>-68.5 0</intersection>
<intersection>-53 9</intersection>
<intersection>-40.5 10</intersection>
<intersection>1 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-112,-68.5,-112</points>
<connection>
<GID>627</GID>
<name>OUT_3</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>1,-159,1,-51.5</points>
<intersection>-159 1</intersection>
<intersection>-51.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>1,-51.5,49,-51.5</points>
<connection>
<GID>613</GID>
<name>IN_3</name></connection>
<intersection>1 6</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-53,-159,-53,-107</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-40.5,-159,-40.5,-107</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection></vsegment></shape></wire>
<wire>
<ID>961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,-160.5,-69,-113</points>
<intersection>-160.5 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-160.5,2,-160.5</points>
<intersection>-69 0</intersection>
<intersection>-53 4</intersection>
<intersection>-40.5 5</intersection>
<intersection>2 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-113,-69,-113</points>
<connection>
<GID>627</GID>
<name>OUT_2</name></connection>
<intersection>-69 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2,-160.5,2,-52.5</points>
<intersection>-160.5 1</intersection>
<intersection>-52.5 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-53,-160.5,-53,-118</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-40.5,-160.5,-40.5,-118</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>2,-52.5,49,-52.5</points>
<connection>
<GID>613</GID>
<name>IN_2</name></connection>
<intersection>2 3</intersection></hsegment></shape></wire>
<wire>
<ID>962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,-161.5,-69.5,-114</points>
<intersection>-161.5 1</intersection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,-161.5,3,-161.5</points>
<intersection>-69.5 0</intersection>
<intersection>-53 8</intersection>
<intersection>-40.5 9</intersection>
<intersection>3 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-114,-69.5,-114</points>
<connection>
<GID>627</GID>
<name>OUT_1</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>3,-161.5,3,-53.5</points>
<intersection>-161.5 1</intersection>
<intersection>-53.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>3,-53.5,49,-53.5</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<intersection>3 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-53,-161.5,-53,-128.5</points>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>-161.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-40.5,-161.5,-40.5,-128.5</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-161.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-90.5,-28.5,-61.5</points>
<intersection>-90.5 2</intersection>
<intersection>-80 3</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-61.5,-28.5,-61.5</points>
<connection>
<GID>628</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-90.5,-16.5,-90.5</points>
<connection>
<GID>636</GID>
<name>IN_7</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,-80,4.5,-80</points>
<connection>
<GID>668</GID>
<name>IN_7</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>964</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-91.5,-28.5,-72.5</points>
<intersection>-91.5 2</intersection>
<intersection>-81 4</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-72.5,-28.5,-72.5</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-91.5,-16.5,-91.5</points>
<connection>
<GID>636</GID>
<name>IN_6</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-28.5,-81,4.5,-81</points>
<connection>
<GID>668</GID>
<name>IN_6</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>965</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-92.5,-28.5,-82</points>
<intersection>-92.5 2</intersection>
<intersection>-83.5 1</intersection>
<intersection>-82 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-83.5,-28.5,-83.5</points>
<connection>
<GID>630</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-92.5,-16.5,-92.5</points>
<connection>
<GID>636</GID>
<name>IN_5</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,-82,4.5,-82</points>
<connection>
<GID>668</GID>
<name>IN_5</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>966</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-93.5,-16.5,-93.5</points>
<connection>
<GID>636</GID>
<name>IN_4</name></connection>
<intersection>-47 6</intersection>
<intersection>-27.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-27.5,-93.5,-27.5,-83</points>
<intersection>-93.5 1</intersection>
<intersection>-83 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-27.5,-83,4.5,-83</points>
<connection>
<GID>668</GID>
<name>IN_4</name></connection>
<intersection>-27.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-47,-93.5,-47,-93</points>
<connection>
<GID>631</GID>
<name>OUT</name></connection>
<intersection>-93.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>967</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-104,-28.5,-94.5</points>
<intersection>-104 1</intersection>
<intersection>-94.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-104,-28.5,-104</points>
<connection>
<GID>632</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-94.5,-16.5,-94.5</points>
<connection>
<GID>636</GID>
<name>IN_3</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-26.5,-94.5,-26.5,-84</points>
<intersection>-94.5 2</intersection>
<intersection>-84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-26.5,-84,4.5,-84</points>
<connection>
<GID>668</GID>
<name>IN_3</name></connection>
<intersection>-26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-115,-28.5,-95.5</points>
<intersection>-115 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-115,-28.5,-115</points>
<connection>
<GID>633</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-95.5,-16.5,-95.5</points>
<connection>
<GID>636</GID>
<name>IN_2</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25.5,-95.5,-25.5,-85</points>
<intersection>-95.5 2</intersection>
<intersection>-85 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25.5,-85,4.5,-85</points>
<connection>
<GID>668</GID>
<name>IN_2</name></connection>
<intersection>-25.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>969</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-125.5,-28.5,-96.5</points>
<intersection>-125.5 1</intersection>
<intersection>-96.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-125.5,-28.5,-125.5</points>
<connection>
<GID>634</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,-96.5,-16.5,-96.5</points>
<connection>
<GID>636</GID>
<name>IN_1</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24.5,-96.5,-24.5,-86</points>
<intersection>-96.5 2</intersection>
<intersection>-86 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-24.5,-86,4.5,-86</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<intersection>-24.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>970</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-136.5,-28.5,-97.5</points>
<intersection>-136.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28.5,-97.5,-16.5,-97.5</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>-28.5 0</intersection>
<intersection>-23.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-136.5,-28.5,-136.5</points>
<connection>
<GID>635</GID>
<name>OUT</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-23.5,-97.5,-23.5,-87</points>
<intersection>-97.5 1</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-23.5,-87,4.5,-87</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-23.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>971</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,-163,-70,-115</points>
<intersection>-163 1</intersection>
<intersection>-115 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70,-163,4,-163</points>
<intersection>-70 0</intersection>
<intersection>-53 14</intersection>
<intersection>-40.5 15</intersection>
<intersection>4 13</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,-115,-70,-115</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<intersection>-70 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>4,-163,4,-54.5</points>
<intersection>-163 1</intersection>
<intersection>-54.5 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-53,-163,-53,-139.5</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>-163 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-40.5,-163,-40.5,-139.5</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>-163 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>4,-54.5,49,-54.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>4 13</intersection></hsegment></shape></wire>
<wire>
<ID>972</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-120.5,-80,-77.5</points>
<intersection>-120.5 10</intersection>
<intersection>-117 8</intersection>
<intersection>-104 7</intersection>
<intersection>-90.5 6</intersection>
<intersection>-77.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-80,-77.5,-76.5,-77.5</points>
<connection>
<GID>202</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-80,-90.5,-76.5,-90.5</points>
<connection>
<GID>203</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-80,-104,-76.5,-104</points>
<connection>
<GID>626</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-80,-117,-76.5,-117</points>
<connection>
<GID>627</GID>
<name>clock</name></connection>
<intersection>-80 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-83,-120.5,-80,-120.5</points>
<connection>
<GID>638</GID>
<name>CLK</name></connection>
<intersection>-80 0</intersection></hsegment></shape></wire>
<wire>
<ID>973</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-131.5,-49,-53.5</points>
<connection>
<GID>635</GID>
<name>SEL_0</name></connection>
<connection>
<GID>634</GID>
<name>SEL_0</name></connection>
<connection>
<GID>633</GID>
<name>SEL_0</name></connection>
<connection>
<GID>632</GID>
<name>SEL_0</name></connection>
<connection>
<GID>631</GID>
<name>SEL_0</name></connection>
<connection>
<GID>630</GID>
<name>SEL_0</name></connection>
<connection>
<GID>629</GID>
<name>SEL_0</name></connection>
<connection>
<GID>628</GID>
<name>SEL_0</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-102.5,-53.5,-49,-53.5</points>
<intersection>-102.5 2</intersection>
<intersection>-49 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-102.5,-79.5,-102.5,-53.5</points>
<intersection>-79.5 3</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-79.5,-102.5,-79.5</points>
<connection>
<GID>637</GID>
<name>OUT_0</name></connection>
<intersection>-102.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>974</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-131.5,-50,-54</points>
<connection>
<GID>635</GID>
<name>SEL_1</name></connection>
<connection>
<GID>634</GID>
<name>SEL_1</name></connection>
<connection>
<GID>633</GID>
<name>SEL_1</name></connection>
<connection>
<GID>632</GID>
<name>SEL_1</name></connection>
<connection>
<GID>631</GID>
<name>SEL_1</name></connection>
<connection>
<GID>630</GID>
<name>SEL_1</name></connection>
<connection>
<GID>629</GID>
<name>SEL_1</name></connection>
<connection>
<GID>628</GID>
<name>SEL_1</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,-54,-50,-54</points>
<intersection>-103 2</intersection>
<intersection>-50 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-103,-77.5,-103,-54</points>
<intersection>-77.5 3</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-77.5,-103,-77.5</points>
<connection>
<GID>637</GID>
<name>OUT_1</name></connection>
<intersection>-103 2</intersection></hsegment></shape></wire>
<wire>
<ID>975</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-101,-34,-61.5</points>
<intersection>-101 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-61.5,-34,-61.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-101,-14.5,-101</points>
<connection>
<GID>653</GID>
<name>IN_7</name></connection>
<intersection>-34 0</intersection>
<intersection>-28 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-28,-111.5,-28,-101</points>
<intersection>-111.5 4</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-28,-111.5,4.5,-111.5</points>
<connection>
<GID>670</GID>
<name>IN_7</name></connection>
<intersection>-28 3</intersection></hsegment></shape></wire>
<wire>
<ID>976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-102,-34,-72.5</points>
<intersection>-102 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-72.5,-34,-72.5</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-102,-14.5,-102</points>
<connection>
<GID>653</GID>
<name>IN_6</name></connection>
<intersection>-34 0</intersection>
<intersection>-27.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-112.5,-27.5,-102</points>
<intersection>-112.5 4</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-27.5,-112.5,4.5,-112.5</points>
<connection>
<GID>670</GID>
<name>IN_6</name></connection>
<intersection>-27.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-103,-34,-83.5</points>
<intersection>-103 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-83.5,-34,-83.5</points>
<connection>
<GID>647</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-103,-14.5,-103</points>
<connection>
<GID>653</GID>
<name>IN_5</name></connection>
<intersection>-34 0</intersection>
<intersection>-25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25.5,-113.5,-25.5,-103</points>
<intersection>-113.5 4</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25.5,-113.5,4.5,-113.5</points>
<connection>
<GID>670</GID>
<name>IN_5</name></connection>
<intersection>-25.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-104,-34,-93</points>
<intersection>-104 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-93,-34,-93</points>
<connection>
<GID>648</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-104,-14.5,-104</points>
<connection>
<GID>653</GID>
<name>IN_4</name></connection>
<intersection>-34 0</intersection>
<intersection>-24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24,-114.5,-24,-104</points>
<intersection>-114.5 4</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-24,-114.5,4.5,-114.5</points>
<connection>
<GID>670</GID>
<name>IN_4</name></connection>
<intersection>-24 3</intersection></hsegment></shape></wire>
<wire>
<ID>979</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-34,-105,-14.5,-105</points>
<connection>
<GID>653</GID>
<name>IN_3</name></connection>
<intersection>-34 2</intersection>
<intersection>-22 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34,-105,-34,-104</points>
<intersection>-105 1</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-34.5,-104,-34,-104</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>-34 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22,-115.5,-22,-105</points>
<intersection>-115.5 5</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-22,-115.5,4.5,-115.5</points>
<connection>
<GID>670</GID>
<name>IN_3</name></connection>
<intersection>-22 4</intersection></hsegment></shape></wire>
<wire>
<ID>980</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-115,-34,-106</points>
<intersection>-115 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-115,-34,-115</points>
<connection>
<GID>650</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-106,-14.5,-106</points>
<connection>
<GID>653</GID>
<name>IN_2</name></connection>
<intersection>-34 0</intersection>
<intersection>-20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-20,-116.5,-20,-106</points>
<intersection>-116.5 4</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20,-116.5,4.5,-116.5</points>
<connection>
<GID>670</GID>
<name>IN_2</name></connection>
<intersection>-20 3</intersection></hsegment></shape></wire>
<wire>
<ID>981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-125.5,-34,-107</points>
<intersection>-125.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-125.5,-34,-125.5</points>
<connection>
<GID>651</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34,-107,-14.5,-107</points>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<intersection>-34 0</intersection>
<intersection>-19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19,-117.5,-19,-107</points>
<intersection>-117.5 4</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-19,-117.5,4.5,-117.5</points>
<connection>
<GID>670</GID>
<name>IN_1</name></connection>
<intersection>-19 3</intersection></hsegment></shape></wire>
<wire>
<ID>982</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-136.5,-34,-108</points>
<intersection>-136.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-108,-14.5,-108</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection>
<intersection>-18 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,-136.5,-34,-136.5</points>
<connection>
<GID>652</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,-118.5,-18,-108</points>
<intersection>-118.5 4</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-18,-118.5,4.5,-118.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>983</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,-131.5,-36.5,-55</points>
<connection>
<GID>652</GID>
<name>SEL_0</name></connection>
<connection>
<GID>651</GID>
<name>SEL_0</name></connection>
<connection>
<GID>650</GID>
<name>SEL_0</name></connection>
<connection>
<GID>649</GID>
<name>SEL_0</name></connection>
<connection>
<GID>648</GID>
<name>SEL_0</name></connection>
<connection>
<GID>647</GID>
<name>SEL_0</name></connection>
<connection>
<GID>646</GID>
<name>SEL_0</name></connection>
<connection>
<GID>645</GID>
<name>SEL_0</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-101.5,-55,-36.5,-55</points>
<intersection>-101.5 2</intersection>
<intersection>-36.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-101.5,-93.5,-101.5,-55</points>
<intersection>-93.5 3</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-93.5,-101.5,-93.5</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-131.5,-37.5,-54.5</points>
<connection>
<GID>652</GID>
<name>SEL_1</name></connection>
<connection>
<GID>651</GID>
<name>SEL_1</name></connection>
<connection>
<GID>650</GID>
<name>SEL_1</name></connection>
<connection>
<GID>649</GID>
<name>SEL_1</name></connection>
<connection>
<GID>648</GID>
<name>SEL_1</name></connection>
<connection>
<GID>647</GID>
<name>SEL_1</name></connection>
<connection>
<GID>646</GID>
<name>SEL_1</name></connection>
<connection>
<GID>645</GID>
<name>SEL_1</name></connection>
<intersection>-54.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-102,-54.5,-37.5,-54.5</points>
<intersection>-102 16</intersection>
<intersection>-37.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-102,-91.5,-102,-54.5</points>
<intersection>-91.5 18</intersection>
<intersection>-54.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-103.5,-91.5,-102,-91.5</points>
<connection>
<GID>644</GID>
<name>OUT_1</name></connection>
<intersection>-102 16</intersection></hsegment></shape></wire>
<wire>
<ID>985</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-108,-81,-68.5</points>
<intersection>-108 6</intersection>
<intersection>-95 3</intersection>
<intersection>-87 4</intersection>
<intersection>-81.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81,-68.5,-79.5,-68.5</points>
<connection>
<GID>202</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-81,-81.5,-79.5,-81.5</points>
<connection>
<GID>203</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-81,-95,-79.5,-95</points>
<connection>
<GID>626</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-87.5,-87,-81,-87</points>
<connection>
<GID>655</GID>
<name>OUT_3</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-81,-108,-79.5,-108</points>
<connection>
<GID>627</GID>
<name>IN_7</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>986</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,-109,-81.5,-69.5</points>
<intersection>-109 6</intersection>
<intersection>-96 5</intersection>
<intersection>-89 2</intersection>
<intersection>-82.5 3</intersection>
<intersection>-69.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-89,-81.5,-89</points>
<connection>
<GID>655</GID>
<name>OUT_2</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-81.5,-82.5,-79.5,-82.5</points>
<connection>
<GID>203</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-81.5,-69.5,-79.5,-69.5</points>
<connection>
<GID>202</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-81.5,-96,-79.5,-96</points>
<connection>
<GID>626</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-81.5,-109,-79.5,-109</points>
<connection>
<GID>627</GID>
<name>IN_6</name></connection>
<intersection>-81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82,-110,-82,-70.5</points>
<intersection>-110 6</intersection>
<intersection>-97 3</intersection>
<intersection>-91 2</intersection>
<intersection>-83.5 4</intersection>
<intersection>-70.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-91,-82,-91</points>
<connection>
<GID>655</GID>
<name>OUT_1</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-82,-97,-79.5,-97</points>
<connection>
<GID>626</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-82,-83.5,-79.5,-83.5</points>
<connection>
<GID>203</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-82,-70.5,-79.5,-70.5</points>
<connection>
<GID>202</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-82,-110,-79.5,-110</points>
<connection>
<GID>627</GID>
<name>IN_5</name></connection>
<intersection>-82 0</intersection></hsegment></shape></wire>
<wire>
<ID>988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82.5,-111,-82.5,-71.5</points>
<intersection>-111 6</intersection>
<intersection>-98 3</intersection>
<intersection>-93 2</intersection>
<intersection>-84.5 4</intersection>
<intersection>-71.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-93,-82.5,-93</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-82.5,-98,-79.5,-98</points>
<connection>
<GID>626</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-82.5,-84.5,-79.5,-84.5</points>
<connection>
<GID>203</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-82.5,-71.5,-79.5,-71.5</points>
<connection>
<GID>202</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-82.5,-111,-79.5,-111</points>
<connection>
<GID>627</GID>
<name>IN_4</name></connection>
<intersection>-82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83,-112,-83,-72.5</points>
<intersection>-112 5</intersection>
<intersection>-99 2</intersection>
<intersection>-85.5 3</intersection>
<intersection>-72.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-99,-79.5,-99</points>
<connection>
<GID>626</GID>
<name>IN_3</name></connection>
<connection>
<GID>656</GID>
<name>OUT_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-83,-85.5,-79.5,-85.5</points>
<connection>
<GID>203</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-83,-72.5,-79.5,-72.5</points>
<connection>
<GID>202</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-83,-112,-79.5,-112</points>
<connection>
<GID>627</GID>
<name>IN_3</name></connection>
<intersection>-83 0</intersection></hsegment></shape></wire>
<wire>
<ID>990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83.5,-113,-83.5,-73.5</points>
<intersection>-113 5</intersection>
<intersection>-101 2</intersection>
<intersection>-100 4</intersection>
<intersection>-86.5 3</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83.5,-73.5,-79.5,-73.5</points>
<connection>
<GID>202</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-101,-83.5,-101</points>
<connection>
<GID>656</GID>
<name>OUT_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-83.5,-86.5,-79.5,-86.5</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-83.5,-100,-79.5,-100</points>
<connection>
<GID>626</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-83.5,-113,-79.5,-113</points>
<connection>
<GID>627</GID>
<name>IN_2</name></connection>
<intersection>-83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84,-114,-84,-74.5</points>
<intersection>-114 5</intersection>
<intersection>-103 2</intersection>
<intersection>-101 4</intersection>
<intersection>-87.5 3</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84,-74.5,-79.5,-74.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-103,-84,-103</points>
<connection>
<GID>656</GID>
<name>OUT_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84,-87.5,-79.5,-87.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84,-101,-79.5,-101</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-84,-114,-79.5,-114</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<intersection>-84 0</intersection></hsegment></shape></wire>
<wire>
<ID>992</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-84.5,-115,-84.5,-75.5</points>
<intersection>-115 5</intersection>
<intersection>-105 2</intersection>
<intersection>-102 4</intersection>
<intersection>-88.5 3</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-84.5,-75.5,-79.5,-75.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,-105,-84.5,-105</points>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-84.5,-88.5,-79.5,-88.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-84.5,-102,-79.5,-102</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-84.5,-115,-79.5,-115</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>-84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>993</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-66.5,-77.5,-58.5</points>
<intersection>-66.5 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-58.5,-77.5,-58.5</points>
<connection>
<GID>658</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-66.5,-76.5,-66.5</points>
<connection>
<GID>202</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>994</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-79.5,-77.5,-57.5</points>
<intersection>-79.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-57.5,-77.5,-57.5</points>
<connection>
<GID>658</GID>
<name>OUT_1</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-79.5,-76.5,-79.5</points>
<connection>
<GID>203</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-93,-77.5,-56.5</points>
<intersection>-93 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-56.5,-77.5,-56.5</points>
<connection>
<GID>658</GID>
<name>OUT_2</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-93,-76.5,-93</points>
<connection>
<GID>626</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>996</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-106,-77.5,-55.5</points>
<intersection>-106 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,-55.5,-77.5,-55.5</points>
<connection>
<GID>658</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-106,-76.5,-106</points>
<connection>
<GID>627</GID>
<name>load</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94.5,-56.5,-93.5,-56.5</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>-93.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-93.5,-56.5,-93.5,-55.5</points>
<connection>
<GID>658</GID>
<name>ENABLE</name></connection>
<intersection>-56.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>998</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89,-72.5,-89,-61.5</points>
<intersection>-72.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94,-61.5,-89,-61.5</points>
<intersection>-94 3</intersection>
<intersection>-89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,-72.5,-89,-72.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>-89 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-94,-61.5,-94,-58.5</points>
<intersection>-61.5 1</intersection>
<intersection>-58.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-94,-58.5,-93.5,-58.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-94 3</intersection></hsegment></shape></wire>
<wire>
<ID>999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,-70.5,-88.5,-61</points>
<intersection>-70.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-61,-88.5,-61</points>
<intersection>-93.5 3</intersection>
<intersection>-88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90.5,-70.5,-88.5,-70.5</points>
<connection>
<GID>661</GID>
<name>OUT_1</name></connection>
<intersection>-88.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-93.5,-61,-93.5,-57.5</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>1000</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-78.5,6.5,-72.5</points>
<connection>
<GID>668</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>672</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-110,6.5,-101</points>
<connection>
<GID>670</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>678</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1004</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-118.5,30.5,-93</points>
<intersection>-118.5 1</intersection>
<intersection>-93 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-118.5,44.5,-118.5</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-93,44.5,-93</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-118.5,44.5,-116</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-118.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1005</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-115,30.5,-87</points>
<intersection>-115 1</intersection>
<intersection>-92 3</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-115,44.5,-115</points>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-87,30.5,-87</points>
<connection>
<GID>668</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-92,44.5,-92</points>
<connection>
<GID>621</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1006</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-117.5,30.5,-91</points>
<intersection>-117.5 2</intersection>
<intersection>-114 1</intersection>
<intersection>-91 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-114,44.5,-114</points>
<connection>
<GID>622</GID>
<name>IN_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-117.5,30.5,-117.5</points>
<connection>
<GID>670</GID>
<name>OUT_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-91,44.5,-91</points>
<connection>
<GID>621</GID>
<name>IN_2</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1007</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-113,30.5,-86</points>
<intersection>-113 1</intersection>
<intersection>-90 3</intersection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-113,44.5,-113</points>
<connection>
<GID>622</GID>
<name>IN_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-86,30.5,-86</points>
<connection>
<GID>668</GID>
<name>OUT_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-90,44.5,-90</points>
<connection>
<GID>621</GID>
<name>IN_3</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1008</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-116.5,30.5,-112</points>
<intersection>-116.5 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-112,44.5,-112</points>
<connection>
<GID>622</GID>
<name>IN_4</name></connection>
<intersection>30.5 0</intersection>
<intersection>39.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-116.5,30.5,-116.5</points>
<connection>
<GID>670</GID>
<name>OUT_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-112,39.5,-89</points>
<intersection>-112 1</intersection>
<intersection>-89 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39.5,-89,44.5,-89</points>
<connection>
<GID>621</GID>
<name>IN_4</name></connection>
<intersection>39.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1009</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-115.5,30.5,-110</points>
<intersection>-115.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-110,44.5,-110</points>
<connection>
<GID>622</GID>
<name>IN_6</name></connection>
<intersection>30.5 0</intersection>
<intersection>44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-115.5,30.5,-115.5</points>
<connection>
<GID>670</GID>
<name>OUT_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-110,44,-87</points>
<intersection>-110 1</intersection>
<intersection>-87 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>44,-87,44.5,-87</points>
<connection>
<GID>621</GID>
<name>IN_6</name></connection>
<intersection>44 3</intersection></hsegment></shape></wire>
<wire>
<ID>1010</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-114.5,30.5,-108</points>
<intersection>-114.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-108,44.5,-108</points>
<connection>
<GID>622</GID>
<name>IN_8</name></connection>
<intersection>30.5 0</intersection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-114.5,30.5,-114.5</points>
<connection>
<GID>670</GID>
<name>OUT_4</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-108,42.5,-83</points>
<intersection>-108 1</intersection>
<intersection>-85 6</intersection>
<intersection>-83 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-83,44.5,-83</points>
<connection>
<GID>621</GID>
<name>IN_10</name></connection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>42.5,-85,44.5,-85</points>
<connection>
<GID>621</GID>
<name>IN_8</name></connection>
<intersection>42.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1011</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-113.5,30.5,-106</points>
<intersection>-113.5 2</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-106,44.5,-106</points>
<connection>
<GID>622</GID>
<name>IN_10</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-113.5,30.5,-113.5</points>
<connection>
<GID>670</GID>
<name>OUT_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1012</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-112.5,30.5,-104</points>
<intersection>-112.5 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-104,44.5,-104</points>
<connection>
<GID>622</GID>
<name>IN_12</name></connection>
<intersection>30.5 0</intersection>
<intersection>43.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-112.5,30.5,-112.5</points>
<connection>
<GID>670</GID>
<name>OUT_6</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-104,43.5,-81</points>
<intersection>-104 1</intersection>
<intersection>-81 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-81,44.5,-81</points>
<connection>
<GID>621</GID>
<name>IN_12</name></connection>
<intersection>43.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1013</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-111.5,30.5,-102</points>
<intersection>-111.5 2</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-102,44.5,-102</points>
<connection>
<GID>622</GID>
<name>IN_14</name></connection>
<intersection>30.5 0</intersection>
<intersection>38 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-111.5,30.5,-111.5</points>
<connection>
<GID>670</GID>
<name>OUT_7</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-102,38,-79</points>
<intersection>-102 1</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,-79,44.5,-79</points>
<connection>
<GID>621</GID>
<name>IN_14</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>1014</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-111,30.5,-85</points>
<intersection>-111 1</intersection>
<intersection>-88 3</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-111,44.5,-111</points>
<connection>
<GID>622</GID>
<name>IN_5</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-85,30.5,-85</points>
<connection>
<GID>668</GID>
<name>OUT_2</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-88,44.5,-88</points>
<connection>
<GID>621</GID>
<name>IN_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-109,30.5,-84</points>
<intersection>-109 1</intersection>
<intersection>-86 3</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-109,44.5,-109</points>
<connection>
<GID>622</GID>
<name>IN_7</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-84,30.5,-84</points>
<connection>
<GID>668</GID>
<name>OUT_3</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-86,44.5,-86</points>
<connection>
<GID>621</GID>
<name>IN_7</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-107,30.5,-83</points>
<intersection>-107 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-107,44.5,-107</points>
<connection>
<GID>622</GID>
<name>IN_9</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-83,44.5,-83</points>
<connection>
<GID>668</GID>
<name>OUT_4</name></connection>
<intersection>30.5 0</intersection>
<intersection>44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44.5,-84,44.5,-83</points>
<connection>
<GID>621</GID>
<name>IN_9</name></connection>
<intersection>-83 2</intersection></vsegment></shape></wire>
<wire>
<ID>1017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-105,30.5,-82</points>
<intersection>-105 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-105,44.5,-105</points>
<connection>
<GID>622</GID>
<name>IN_11</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-82,44.5,-82</points>
<connection>
<GID>621</GID>
<name>IN_11</name></connection>
<connection>
<GID>668</GID>
<name>OUT_5</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-103,30.5,-80</points>
<intersection>-103 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-103,44.5,-103</points>
<connection>
<GID>622</GID>
<name>IN_13</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-80,44.5,-80</points>
<connection>
<GID>621</GID>
<name>IN_13</name></connection>
<intersection>17 4</intersection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17,-81,17,-80</points>
<intersection>-81 5</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>8.5,-81,17,-81</points>
<connection>
<GID>668</GID>
<name>OUT_6</name></connection>
<intersection>17 4</intersection></hsegment></shape></wire>
<wire>
<ID>1019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-101,30.5,-78</points>
<intersection>-101 1</intersection>
<intersection>-79 2</intersection>
<intersection>-78 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-101,44.5,-101</points>
<connection>
<GID>622</GID>
<name>IN_15</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-79,30.5,-79</points>
<intersection>8.5 4</intersection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-78,44.5,-78</points>
<connection>
<GID>621</GID>
<name>IN_15</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-80,8.5,-79</points>
<connection>
<GID>668</GID>
<name>OUT_7</name></connection>
<intersection>-79 2</intersection></vsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-22,18,-16</points>
<intersection>-22 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-16,23.5,-16</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-22,18,-22</points>
<connection>
<GID>592</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-20,18,-15</points>
<intersection>-20 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-15,23.5,-15</points>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-20,18,-20</points>
<connection>
<GID>592</GID>
<name>OUT_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-18,18,-14</points>
<intersection>-18 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-14,23.5,-14</points>
<connection>
<GID>587</GID>
<name>IN_2</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-18,18,-18</points>
<connection>
<GID>592</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-16,18,-13</points>
<intersection>-16 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-13,23.5,-13</points>
<connection>
<GID>587</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-16,18,-16</points>
<connection>
<GID>592</GID>
<name>OUT_3</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-12,18,-10</points>
<intersection>-12 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-12,23.5,-12</points>
<connection>
<GID>587</GID>
<name>IN_4</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-10,18,-10</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-11,18,-8</points>
<intersection>-11 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-11,23.5,-11</points>
<connection>
<GID>587</GID>
<name>IN_5</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-8,18,-8</points>
<connection>
<GID>593</GID>
<name>OUT_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-10,18,-6</points>
<intersection>-10 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-10,23.5,-10</points>
<connection>
<GID>587</GID>
<name>IN_6</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-6,18,-6</points>
<connection>
<GID>593</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-9,23.5,-9</points>
<connection>
<GID>587</GID>
<name>IN_7</name></connection>
<intersection>13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-9,13,-4</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-9,40.5,-9</points>
<connection>
<GID>587</GID>
<name>OUT_7</name></connection>
<connection>
<GID>588</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-10,40.5,-10</points>
<connection>
<GID>587</GID>
<name>OUT_6</name></connection>
<connection>
<GID>588</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-11,40.5,-11</points>
<connection>
<GID>587</GID>
<name>OUT_5</name></connection>
<connection>
<GID>588</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-12,40.5,-12</points>
<connection>
<GID>587</GID>
<name>OUT_4</name></connection>
<connection>
<GID>588</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-13,40.5,-13</points>
<connection>
<GID>587</GID>
<name>OUT_3</name></connection>
<connection>
<GID>588</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-14,40.5,-14</points>
<connection>
<GID>587</GID>
<name>OUT_2</name></connection>
<connection>
<GID>588</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-15,40.5,-15</points>
<connection>
<GID>587</GID>
<name>OUT_1</name></connection>
<connection>
<GID>588</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-16,40.5,-16</points>
<connection>
<GID>587</GID>
<name>OUT_0</name></connection>
<connection>
<GID>588</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-9,54.5,-9</points>
<connection>
<GID>588</GID>
<name>OUT_7</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-10,54.5,-10</points>
<connection>
<GID>588</GID>
<name>OUT_6</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-11,54.5,-11</points>
<connection>
<GID>588</GID>
<name>OUT_5</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-12,54.5,-12</points>
<connection>
<GID>588</GID>
<name>OUT_4</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-13,54.5,-13</points>
<connection>
<GID>588</GID>
<name>OUT_3</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-14,54.5,-14</points>
<connection>
<GID>588</GID>
<name>OUT_2</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-7,43.5,3.5</points>
<connection>
<GID>588</GID>
<name>load</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,3.5,43.5,3.5</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-7,27.5,6</points>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection>
<connection>
<GID>587</GID>
<name>count_enable</name></connection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-6,28.5,-6</points>
<intersection>27.5 0</intersection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-7,28.5,-6</points>
<connection>
<GID>587</GID>
<name>count_up</name></connection>
<intersection>-6 2</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>81.5,-59.5,81.5,-45.5</points>
<connection>
<GID>601</GID>
<name>OUT_0</name></connection>
<connection>
<GID>589</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-15,54.5,-15</points>
<connection>
<GID>588</GID>
<name>OUT_1</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-16,54.5,-16</points>
<connection>
<GID>588</GID>
<name>OUT_0</name></connection>
<connection>
<GID>590</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-47.5,96,-47.5</points>
<connection>
<GID>589</GID>
<name>OUT_7</name></connection>
<connection>
<GID>591</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-48.5,96,-48.5</points>
<connection>
<GID>589</GID>
<name>OUT_6</name></connection>
<connection>
<GID>591</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-49.5,96,-49.5</points>
<connection>
<GID>589</GID>
<name>OUT_5</name></connection>
<connection>
<GID>591</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-50.5,96,-50.5</points>
<connection>
<GID>589</GID>
<name>OUT_4</name></connection>
<connection>
<GID>591</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-51.5,96,-51.5</points>
<connection>
<GID>589</GID>
<name>OUT_3</name></connection>
<connection>
<GID>591</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-52.5,96,-52.5</points>
<connection>
<GID>589</GID>
<name>OUT_2</name></connection>
<connection>
<GID>591</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-53.5,96,-53.5</points>
<connection>
<GID>589</GID>
<name>OUT_1</name></connection>
<connection>
<GID>591</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-54.5,96,-54.5</points>
<connection>
<GID>589</GID>
<name>OUT_0</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-59.5,99,-45.5</points>
<connection>
<GID>591</GID>
<name>load</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-59.5,99,-59.5</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-54.5,107.5,-54.5</points>
<connection>
<GID>591</GID>
<name>OUT_0</name></connection>
<connection>
<GID>607</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-53.5,107.5,-53.5</points>
<connection>
<GID>591</GID>
<name>OUT_1</name></connection>
<connection>
<GID>607</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-43.5,43.5,-18</points>
<connection>
<GID>588</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-43.5,99,-43.5</points>
<connection>
<GID>618</GID>
<name>OUT</name></connection>
<intersection>13.5 6</intersection>
<intersection>43.5 0</intersection>
<intersection>81.5 5</intersection>
<intersection>99 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>99,-56.5,99,-43.5</points>
<connection>
<GID>591</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>81.5,-56.5,81.5,-43.5</points>
<connection>
<GID>589</GID>
<name>clock</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>13.5,-43.5,13.5,-25</points>
<intersection>-43.5 1</intersection>
<intersection>-25 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13.5,-25,19.5,-25</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>13.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-41.5,28.5,-18</points>
<connection>
<GID>599</GID>
<name>OUT_0</name></connection>
<connection>
<GID>587</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-41.5,101,-41.5</points>
<intersection>28.5 0</intersection>
<intersection>45.5 3</intersection>
<intersection>83.5 7</intersection>
<intersection>101 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-41.5,45.5,-18</points>
<connection>
<GID>588</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>101,-56.5,101,-41.5</points>
<connection>
<GID>591</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>83.5,-56.5,83.5,-41.5</points>
<connection>
<GID>589</GID>
<name>clear</name></connection>
<intersection>-41.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-10,67.5,-10</points>
<connection>
<GID>608</GID>
<name>OUT_0</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-25,65.5,-10</points>
<intersection>-25 4</intersection>
<intersection>-12 7</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-25,65.5,-25</points>
<intersection>51 8</intersection>
<intersection>65.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>64.5,-12,65.5,-12</points>
<connection>
<GID>590</GID>
<name>write_enable</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>51,-46,51,-25</points>
<connection>
<GID>613</GID>
<name>ENABLE_0</name></connection>
<intersection>-25 4</intersection></vsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-13,67.5,-13</points>
<connection>
<GID>590</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>609</GID>
<name>OUT_0</name></connection>
<intersection>67.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>67.5,-25,67.5,-13</points>
<intersection>-25 6</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>67.5,-25,73,-25</points>
<intersection>67.5 5</intersection>
<intersection>73 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>73,-46,73,-25</points>
<connection>
<GID>612</GID>
<name>ENABLE_0</name></connection>
<intersection>-25 6</intersection></vsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-53.5,71,-53.5</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<connection>
<GID>613</GID>
<name>OUT_1</name></connection>
<intersection>62 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>62,-53.5,62,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-52.5,71,-52.5</points>
<connection>
<GID>612</GID>
<name>IN_2</name></connection>
<connection>
<GID>613</GID>
<name>OUT_2</name></connection>
<intersection>61 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>61,-52.5,61,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_2</name></connection>
<intersection>-52.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-51.5,71,-51.5</points>
<connection>
<GID>612</GID>
<name>IN_3</name></connection>
<connection>
<GID>613</GID>
<name>OUT_3</name></connection>
<intersection>60 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>60,-51.5,60,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_3</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-50.5,71,-50.5</points>
<connection>
<GID>612</GID>
<name>IN_4</name></connection>
<connection>
<GID>613</GID>
<name>OUT_4</name></connection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-50.5,59,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_4</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-49.5,71,-49.5</points>
<connection>
<GID>612</GID>
<name>IN_5</name></connection>
<connection>
<GID>613</GID>
<name>OUT_5</name></connection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-49.5,58,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_5</name></connection>
<intersection>-49.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-48.5,71,-48.5</points>
<connection>
<GID>612</GID>
<name>IN_6</name></connection>
<connection>
<GID>613</GID>
<name>OUT_6</name></connection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-48.5,57,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_6</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-47.5,71,-47.5</points>
<connection>
<GID>612</GID>
<name>IN_7</name></connection>
<connection>
<GID>613</GID>
<name>OUT_7</name></connection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-47.5,56,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_7</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-49.5,78.5,-49.5</points>
<connection>
<GID>589</GID>
<name>IN_5</name></connection>
<connection>
<GID>612</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-54.5,78.5,-54.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-53.5,78.5,-53.5</points>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<connection>
<GID>612</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-52.5,78.5,-52.5</points>
<connection>
<GID>589</GID>
<name>IN_2</name></connection>
<connection>
<GID>612</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-51.5,78.5,-51.5</points>
<connection>
<GID>589</GID>
<name>IN_3</name></connection>
<connection>
<GID>612</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-50.5,78.5,-50.5</points>
<connection>
<GID>589</GID>
<name>IN_4</name></connection>
<connection>
<GID>612</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-47.5,78.5,-47.5</points>
<connection>
<GID>589</GID>
<name>IN_7</name></connection>
<connection>
<GID>612</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-48.5,78.5,-48.5</points>
<connection>
<GID>589</GID>
<name>IN_6</name></connection>
<connection>
<GID>612</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-54.5,71,-54.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-54.5,63,-19.5</points>
<connection>
<GID>590</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>590</GID>
<name>DATA_IN_0</name></connection>
<intersection>-54.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117.5,-51.5,119.5,-51.5</points>
<connection>
<GID>607</GID>
<name>ENABLE_0</name></connection>
<intersection>119.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>119.5,-51.5,119.5,-30.5</points>
<connection>
<GID>615</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-44.5,5,-44.5</points>
<connection>
<GID>594</GID>
<name>CLK</name></connection>
<connection>
<GID>618</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-42.5,5,-40.5</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-40.5,5,-40.5</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-26,26.5,-18</points>
<connection>
<GID>587</GID>
<name>clock</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-26,26.5,-26</points>
<connection>
<GID>617</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,-27,19.5,-27</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>-1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-27,-1.5,-24.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-7,26.5,1</points>
<connection>
<GID>587</GID>
<name>load</name></connection>
<intersection>1 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-1.5,-18.5,-1.5,1</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,1,26.5,1</points>
<intersection>-1.5 1</intersection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-67.5,35,-67.5</points>
<connection>
<GID>492</GID>
<name>ENABLE</name></connection>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-62,86.5,-62</points>
<intersection>30.5 8</intersection>
<intersection>86.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>86.5,-113.5,86.5,-62</points>
<intersection>-113.5 18</intersection>
<intersection>-108.5 19</intersection>
<intersection>-103.5 20</intersection>
<intersection>-98.5 21</intersection>
<intersection>-93.5 22</intersection>
<intersection>-88.5 23</intersection>
<intersection>-83.5 24</intersection>
<intersection>-78.5 25</intersection>
<intersection>-62 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>30.5,-70.5,30.5,-62</points>
<intersection>-70.5 10</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>30.5,-70.5,35,-70.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>30.5 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>86.5,-113.5,89.5,-113.5</points>
<connection>
<GID>520</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>86.5,-108.5,89.5,-108.5</points>
<connection>
<GID>519</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>86.5,-103.5,89.5,-103.5</points>
<connection>
<GID>518</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>86.5,-98.5,89.5,-98.5</points>
<connection>
<GID>517</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>86.5,-93.5,89.5,-93.5</points>
<connection>
<GID>516</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>86.5,-88.5,89.5,-88.5</points>
<connection>
<GID>515</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>86.5,-83.5,89.5,-83.5</points>
<connection>
<GID>514</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>86.5,-78.5,89.5,-78.5</points>
<connection>
<GID>513</GID>
<name>SEL_0</name></connection>
<intersection>86.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-99.5,42,-70.5</points>
<intersection>-99.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-70.5,42,-70.5</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-99.5,46.5,-99.5</points>
<connection>
<GID>622</GID>
<name>ENABLE_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-76.5,46.5,-69.5</points>
<connection>
<GID>621</GID>
<name>ENABLE_0</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-69.5,46.5,-69.5</points>
<connection>
<GID>492</GID>
<name>OUT_1</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-112.5,63,-112.5</points>
<connection>
<GID>497</GID>
<name>carry_out</name></connection>
<connection>
<GID>498</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-116,50,-99.5</points>
<intersection>-116 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-99.5,60,-99.5</points>
<connection>
<GID>497</GID>
<name>IN_B_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-116,50,-116</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-114,50.5,-100.5</points>
<intersection>-114 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-100.5,60,-100.5</points>
<connection>
<GID>497</GID>
<name>IN_B_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-114,50.5,-114</points>
<connection>
<GID>622</GID>
<name>OUT_2</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-112,51,-101.5</points>
<intersection>-112 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-101.5,60,-101.5</points>
<connection>
<GID>497</GID>
<name>IN_B_2</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-112,51,-112</points>
<connection>
<GID>622</GID>
<name>OUT_4</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-110,51.5,-102.5</points>
<intersection>-110 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-102.5,60,-102.5</points>
<connection>
<GID>497</GID>
<name>IN_B_3</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-110,51.5,-110</points>
<connection>
<GID>622</GID>
<name>OUT_6</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>395.224,21.0892,786.705,-185.661</PageViewport>
<gate>
<ID>778</ID>
<type>AA_LABEL</type>
<position>662,-142.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>779</ID>
<type>AA_LABEL</type>
<position>647.5,-115</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>780</ID>
<type>AA_LABEL</type>
<position>648,-121.5</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>781</ID>
<type>AA_LABEL</type>
<position>647.5,-131</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>782</ID>
<type>AA_LABEL</type>
<position>648.5,-138</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>649.5,-111</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1105 </input>
<output>
<ID>OUT</ID>1129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AA_AND2</type>
<position>654.5,-107.5</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1107 </input>
<output>
<ID>OUT</ID>1130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>785</ID>
<type>AA_AND2</type>
<position>649.5,-104</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1109 </input>
<output>
<ID>OUT</ID>1131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>AA_AND2</type>
<position>654.5,-100.5</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1111 </input>
<output>
<ID>OUT</ID>1132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>787</ID>
<type>AA_AND2</type>
<position>649.5,-97</position>
<input>
<ID>IN_0</ID>1114 </input>
<input>
<ID>IN_1</ID>1113 </input>
<output>
<ID>OUT</ID>1133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>788</ID>
<type>AA_AND2</type>
<position>654.5,-93.5</position>
<input>
<ID>IN_0</ID>1116 </input>
<input>
<ID>IN_1</ID>1115 </input>
<output>
<ID>OUT</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>789</ID>
<type>AA_AND2</type>
<position>649.5,-90</position>
<input>
<ID>IN_0</ID>1118 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>790</ID>
<type>AA_AND2</type>
<position>654.5,-86.5</position>
<input>
<ID>IN_0</ID>1120 </input>
<input>
<ID>IN_1</ID>1119 </input>
<output>
<ID>OUT</ID>1136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>791</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-98</position>
<input>
<ID>IN_0</ID>1128 </input>
<input>
<ID>IN_1</ID>1136 </input>
<output>
<ID>OUT</ID>1144 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>792</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-103</position>
<input>
<ID>IN_0</ID>1127 </input>
<input>
<ID>IN_1</ID>1135 </input>
<output>
<ID>OUT</ID>1143 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>793</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-108</position>
<input>
<ID>IN_0</ID>1126 </input>
<input>
<ID>IN_1</ID>1134 </input>
<output>
<ID>OUT</ID>1142 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-113</position>
<input>
<ID>IN_0</ID>1125 </input>
<input>
<ID>IN_1</ID>1133 </input>
<output>
<ID>OUT</ID>1141 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>795</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-118</position>
<input>
<ID>IN_0</ID>1124 </input>
<input>
<ID>IN_1</ID>1132 </input>
<output>
<ID>OUT</ID>1140 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>796</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-123</position>
<input>
<ID>IN_0</ID>1123 </input>
<input>
<ID>IN_1</ID>1131 </input>
<output>
<ID>OUT</ID>1139 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>797</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-128</position>
<input>
<ID>IN_0</ID>1122 </input>
<input>
<ID>IN_1</ID>1130 </input>
<output>
<ID>OUT</ID>1138 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>798</ID>
<type>AA_MUX_2x1</type>
<position>679.5,-133</position>
<input>
<ID>IN_0</ID>1121 </input>
<input>
<ID>IN_1</ID>1129 </input>
<output>
<ID>OUT</ID>1137 </output>
<input>
<ID>SEL_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>799</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>725,-116</position>
<input>
<ID>IN_0</ID>1137 </input>
<input>
<ID>IN_1</ID>1138 </input>
<input>
<ID>IN_2</ID>1139 </input>
<input>
<ID>IN_3</ID>1140 </input>
<input>
<ID>IN_4</ID>1141 </input>
<input>
<ID>IN_5</ID>1142 </input>
<input>
<ID>IN_6</ID>1143 </input>
<input>
<ID>IN_7</ID>1144 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_LABEL</type>
<position>679.5,-136.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>801</ID>
<type>AA_LABEL</type>
<position>680.5,-94</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>802</ID>
<type>GA_LED</type>
<position>693.5,-125</position>
<input>
<ID>N_in2</ID>1144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>803</ID>
<type>GA_LED</type>
<position>696,-125</position>
<input>
<ID>N_in2</ID>1143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>804</ID>
<type>GA_LED</type>
<position>698.5,-125</position>
<input>
<ID>N_in2</ID>1142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>805</ID>
<type>GA_LED</type>
<position>701,-125</position>
<input>
<ID>N_in2</ID>1141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>806</ID>
<type>GA_LED</type>
<position>703.5,-125</position>
<input>
<ID>N_in2</ID>1140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>807</ID>
<type>GA_LED</type>
<position>706,-125</position>
<input>
<ID>N_in2</ID>1139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>808</ID>
<type>GA_LED</type>
<position>708.5,-125</position>
<input>
<ID>N_in2</ID>1138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>809</ID>
<type>GA_LED</type>
<position>711,-125</position>
<input>
<ID>N_in2</ID>1137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>810</ID>
<type>AA_LABEL</type>
<position>711,-127</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>811</ID>
<type>AA_LABEL</type>
<position>708.5,-127</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>812</ID>
<type>AA_LABEL</type>
<position>706,-127</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>813</ID>
<type>AA_LABEL</type>
<position>703.5,-127</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>814</ID>
<type>AA_LABEL</type>
<position>701,-127</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>815</ID>
<type>AA_LABEL</type>
<position>698.5,-127</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>816</ID>
<type>AA_LABEL</type>
<position>696,-127</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>817</ID>
<type>AA_LABEL</type>
<position>693.5,-127</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>819</ID>
<type>AA_LABEL</type>
<position>483.5,-67.5</position>
<gparam>LABEL_TEXT Control 1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>820</ID>
<type>AA_LABEL</type>
<position>613,-83.5</position>
<gparam>LABEL_TEXT Control 2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>821</ID>
<type>AA_LABEL</type>
<position>623,-82</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>822</ID>
<type>AA_LABEL</type>
<position>563,-41</position>
<gparam>LABEL_TEXT Control 4</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>823</ID>
<type>AA_LABEL</type>
<position>631,-81.5</position>
<gparam>LABEL_TEXT Control 3</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>824</ID>
<type>AA_LABEL</type>
<position>623.5,-9.5</position>
<gparam>LABEL_TEXT Control 5</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>826</ID>
<type>AA_INVERTER</type>
<position>647.5,-45.5</position>
<input>
<ID>IN_0</ID>1060 </input>
<output>
<ID>OUT_0</ID>1232 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>827</ID>
<type>AA_LABEL</type>
<position>655.5,-23</position>
<gparam>LABEL_TEXT Control 6</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>832</ID>
<type>EE_VDD</type>
<position>673.5,-59.5</position>
<output>
<ID>OUT_0</ID>838 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>833</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>621.5,-102.5</position>
<input>
<ID>ENABLE_0</ID>848 </input>
<input>
<ID>IN_0</ID>1257 </input>
<input>
<ID>IN_1</ID>1249 </input>
<input>
<ID>IN_10</ID>1252 </input>
<input>
<ID>IN_11</ID>1245 </input>
<input>
<ID>IN_12</ID>1251 </input>
<input>
<ID>IN_13</ID>1245 </input>
<input>
<ID>IN_14</ID>1250 </input>
<input>
<ID>IN_15</ID>1245 </input>
<input>
<ID>IN_2</ID>1256 </input>
<input>
<ID>IN_3</ID>1248 </input>
<input>
<ID>IN_4</ID>1255 </input>
<input>
<ID>IN_5</ID>1247 </input>
<input>
<ID>IN_6</ID>1254 </input>
<input>
<ID>IN_7</ID>1245 </input>
<input>
<ID>IN_8</ID>1253 </input>
<input>
<ID>IN_9</ID>1245 </input>
<output>
<ID>OUT_0</ID>1330 </output>
<output>
<ID>OUT_1</ID>1323 </output>
<output>
<ID>OUT_10</ID>1335 </output>
<output>
<ID>OUT_11</ID>1336 </output>
<output>
<ID>OUT_12</ID>1333 </output>
<output>
<ID>OUT_13</ID>1331 </output>
<output>
<ID>OUT_14</ID>1334 </output>
<output>
<ID>OUT_15</ID>1338 </output>
<output>
<ID>OUT_2</ID>1327 </output>
<output>
<ID>OUT_3</ID>1326 </output>
<output>
<ID>OUT_4</ID>1324 </output>
<output>
<ID>OUT_5</ID>1325 </output>
<output>
<ID>OUT_6</ID>1328 </output>
<output>
<ID>OUT_7</ID>1329 </output>
<output>
<ID>OUT_8</ID>1337 </output>
<output>
<ID>OUT_9</ID>1332 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>834</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>621.5,-125.5</position>
<input>
<ID>ENABLE_0</ID>847 </input>
<input>
<ID>IN_0</ID>1257 </input>
<input>
<ID>IN_1</ID>1249 </input>
<input>
<ID>IN_10</ID>1252 </input>
<input>
<ID>IN_11</ID>1245 </input>
<input>
<ID>IN_12</ID>1251 </input>
<input>
<ID>IN_13</ID>1245 </input>
<input>
<ID>IN_14</ID>1250 </input>
<input>
<ID>IN_15</ID>1245 </input>
<input>
<ID>IN_2</ID>1256 </input>
<input>
<ID>IN_3</ID>1248 </input>
<input>
<ID>IN_4</ID>1255 </input>
<input>
<ID>IN_5</ID>1247 </input>
<input>
<ID>IN_6</ID>1254 </input>
<input>
<ID>IN_7</ID>1245 </input>
<input>
<ID>IN_8</ID>1253 </input>
<input>
<ID>IN_9</ID>1245 </input>
<output>
<ID>OUT_0</ID>1307 </output>
<output>
<ID>OUT_1</ID>1309 </output>
<output>
<ID>OUT_10</ID>1316 </output>
<output>
<ID>OUT_11</ID>1318 </output>
<output>
<ID>OUT_12</ID>1319 </output>
<output>
<ID>OUT_13</ID>1321 </output>
<output>
<ID>OUT_14</ID>1320 </output>
<output>
<ID>OUT_15</ID>1322 </output>
<output>
<ID>OUT_2</ID>1308 </output>
<output>
<ID>OUT_3</ID>1310 </output>
<output>
<ID>OUT_4</ID>1311 </output>
<output>
<ID>OUT_5</ID>1312 </output>
<output>
<ID>OUT_6</ID>1314 </output>
<output>
<ID>OUT_7</ID>1313 </output>
<output>
<ID>OUT_8</ID>1317 </output>
<output>
<ID>OUT_9</ID>1315 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_OR2</type>
<position>598.5,-89</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_LABEL</type>
<position>602.5,-88.5</position>
<gparam>LABEL_TEXT LD/ST - PC+Off4</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>491</ID>
<type>AA_LABEL</type>
<position>596,-143.5</position>
<gparam>LABEL_TEXT Current PC</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>EE_VDD</type>
<position>581,-93</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>709.5,-57.5</position>
<input>
<ID>IN_0</ID>883 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>831 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>437,-88</position>
<input>
<ID>ENABLE_0</ID>830 </input>
<input>
<ID>IN_0</ID>884 </input>
<output>
<ID>OUT_0</ID>1186 </output>
<output>
<ID>OUT_1</ID>1187 </output>
<output>
<ID>OUT_2</ID>1196 </output>
<output>
<ID>OUT_3</ID>1197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND2</type>
<position>694.5,-65</position>
<input>
<ID>IN_0</ID>833 </input>
<input>
<ID>IN_1</ID>835 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>719.5,-134.5</position>
<input>
<ID>ENABLE_0</ID>196 </input>
<input>
<ID>IN_0</ID>1137 </input>
<input>
<ID>IN_1</ID>1138 </input>
<input>
<ID>IN_2</ID>1139 </input>
<input>
<ID>IN_3</ID>1140 </input>
<input>
<ID>IN_4</ID>1141 </input>
<input>
<ID>IN_5</ID>1142 </input>
<input>
<ID>IN_6</ID>1143 </input>
<input>
<ID>IN_7</ID>1144 </input>
<output>
<ID>OUT_0</ID>270 </output>
<output>
<ID>OUT_1</ID>754 </output>
<output>
<ID>OUT_2</ID>755 </output>
<output>
<ID>OUT_3</ID>756 </output>
<output>
<ID>OUT_4</ID>757 </output>
<output>
<ID>OUT_5</ID>758 </output>
<output>
<ID>OUT_6</ID>759 </output>
<output>
<ID>OUT_7</ID>760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>129</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>437,-108.5</position>
<input>
<ID>ENABLE_0</ID>831 </input>
<input>
<ID>IN_0</ID>883 </input>
<output>
<ID>OUT_0</ID>768 </output>
<output>
<ID>OUT_1</ID>767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>130</ID>
<type>EE_VDD</type>
<position>719.5,-127</position>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND2</type>
<position>694.5,-70.5</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_AND2</type>
<position>694.5,-76</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>835 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>BE_NOR2</type>
<position>687,-61</position>
<input>
<ID>IN_0</ID>761 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>BA_DECODER_2x4</type>
<position>694.5,-57</position>
<input>
<ID>ENABLE</ID>851 </input>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>882 </input>
<output>
<ID>OUT_0</ID>197 </output>
<output>
<ID>OUT_1</ID>883 </output>
<output>
<ID>OUT_2</ID>885 </output>
<output>
<ID>OUT_3</ID>884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>694.5,-53</position>
<gparam>LABEL_TEXT LD/STR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>694,-67.5</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>694,-61.5</position>
<gparam>LABEL_TEXT ADD</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>694,-73</position>
<gparam>LABEL_TEXT BRnzp</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>DM_NOR8</type>
<position>718,-95.5</position>
<input>
<ID>IN_0</ID>1144 </input>
<input>
<ID>IN_1</ID>1143 </input>
<input>
<ID>IN_2</ID>1142 </input>
<input>
<ID>IN_3</ID>1141 </input>
<input>
<ID>IN_4</ID>1137 </input>
<input>
<ID>IN_5</ID>1138 </input>
<input>
<ID>IN_6</ID>1139 </input>
<input>
<ID>IN_7</ID>1140 </input>
<output>
<ID>OUT</ID>762 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>150</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>570,-21</position>
<input>
<ID>ENABLE_0</ID>213 </input>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>215 </input>
<input>
<ID>IN_2</ID>228 </input>
<input>
<ID>IN_3</ID>229 </input>
<input>
<ID>IN_4</ID>230 </input>
<input>
<ID>IN_5</ID>231 </input>
<input>
<ID>IN_6</ID>232 </input>
<input>
<ID>IN_7</ID>233 </input>
<output>
<ID>OUT_0</ID>200 </output>
<output>
<ID>OUT_1</ID>201 </output>
<output>
<ID>OUT_2</ID>204 </output>
<output>
<ID>OUT_3</ID>205 </output>
<output>
<ID>OUT_4</ID>206 </output>
<output>
<ID>OUT_5</ID>207 </output>
<output>
<ID>OUT_6</ID>208 </output>
<output>
<ID>OUT_7</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>540</ID>
<type>AA_LABEL</type>
<position>595.5,-119.5</position>
<gparam>LABEL_TEXT SEXT-Off4</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>541</ID>
<type>AE_SMALL_INVERTER</type>
<position>580.5,-38</position>
<input>
<ID>IN_0</ID>832 </input>
<output>
<ID>OUT_0</ID>849 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>570,-33</position>
<input>
<ID>ENABLE_0</ID>212 </input>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>754 </input>
<input>
<ID>IN_2</ID>755 </input>
<input>
<ID>IN_3</ID>756 </input>
<input>
<ID>IN_4</ID>757 </input>
<input>
<ID>IN_5</ID>758 </input>
<input>
<ID>IN_6</ID>759 </input>
<input>
<ID>IN_7</ID>760 </input>
<output>
<ID>OUT_0</ID>200 </output>
<output>
<ID>OUT_1</ID>201 </output>
<output>
<ID>OUT_2</ID>204 </output>
<output>
<ID>OUT_3</ID>205 </output>
<output>
<ID>OUT_4</ID>206 </output>
<output>
<ID>OUT_5</ID>207 </output>
<output>
<ID>OUT_6</ID>208 </output>
<output>
<ID>OUT_7</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>542</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>597.5,4</position>
<input>
<ID>ENABLE_0</ID>851 </input>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>754 </input>
<input>
<ID>IN_2</ID>755 </input>
<input>
<ID>IN_3</ID>756 </input>
<input>
<ID>IN_4</ID>757 </input>
<input>
<ID>IN_5</ID>758 </input>
<input>
<ID>IN_6</ID>759 </input>
<input>
<ID>IN_7</ID>760 </input>
<output>
<ID>OUT_0</ID>871 </output>
<output>
<ID>OUT_1</ID>872 </output>
<output>
<ID>OUT_2</ID>873 </output>
<output>
<ID>OUT_3</ID>876 </output>
<output>
<ID>OUT_4</ID>875 </output>
<output>
<ID>OUT_5</ID>877 </output>
<output>
<ID>OUT_6</ID>874 </output>
<output>
<ID>OUT_7</ID>878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>155</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>583,-29</position>
<input>
<ID>ENABLE_0</ID>210 </input>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>201 </input>
<input>
<ID>IN_2</ID>204 </input>
<input>
<ID>IN_3</ID>205 </input>
<input>
<ID>IN_4</ID>206 </input>
<input>
<ID>IN_5</ID>207 </input>
<input>
<ID>IN_6</ID>208 </input>
<input>
<ID>IN_7</ID>209 </input>
<output>
<ID>OUT_0</ID>243 </output>
<output>
<ID>OUT_1</ID>249 </output>
<output>
<ID>OUT_2</ID>250 </output>
<output>
<ID>OUT_3</ID>248 </output>
<output>
<ID>OUT_4</ID>263 </output>
<output>
<ID>OUT_5</ID>235 </output>
<output>
<ID>OUT_6</ID>234 </output>
<output>
<ID>OUT_7</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>156</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>595.5,-114.5</position>
<input>
<ID>ENABLE_0</ID>851 </input>
<input>
<ID>IN_3</ID>845 </input>
<input>
<ID>IN_4</ID>843 </input>
<input>
<ID>IN_5</ID>842 </input>
<input>
<ID>IN_6</ID>841 </input>
<output>
<ID>OUT_3</ID>1249 </output>
<output>
<ID>OUT_4</ID>1248 </output>
<output>
<ID>OUT_5</ID>1247 </output>
<output>
<ID>OUT_6</ID>1245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>546</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>607,-9.5</position>
<input>
<ID>ENABLE_0</ID>879 </input>
<input>
<ID>IN_0</ID>867 </input>
<input>
<ID>IN_1</ID>860 </input>
<input>
<ID>IN_2</ID>861 </input>
<input>
<ID>IN_3</ID>864 </input>
<input>
<ID>IN_4</ID>870 </input>
<input>
<ID>IN_5</ID>865 </input>
<input>
<ID>IN_6</ID>866 </input>
<input>
<ID>IN_7</ID>869 </input>
<output>
<ID>OUT_0</ID>871 </output>
<output>
<ID>OUT_1</ID>872 </output>
<output>
<ID>OUT_2</ID>873 </output>
<output>
<ID>OUT_3</ID>876 </output>
<output>
<ID>OUT_4</ID>875 </output>
<output>
<ID>OUT_5</ID>877 </output>
<output>
<ID>OUT_6</ID>874 </output>
<output>
<ID>OUT_7</ID>878 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>547</ID>
<type>AA_TOGGLE</type>
<position>591.5,-43</position>
<output>
<ID>OUT_0</ID>852 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>158</ID>
<type>BA_DECODER_2x4</type>
<position>565,-12</position>
<input>
<ID>ENABLE</ID>210 </input>
<input>
<ID>IN_0</ID>211 </input>
<output>
<ID>OUT_0</ID>212 </output>
<output>
<ID>OUT_1</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>548</ID>
<type>AE_SMALL_INVERTER</type>
<position>607,-2.5</position>
<input>
<ID>IN_0</ID>851 </input>
<output>
<ID>OUT_0</ID>879 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>EE_VDD</type>
<position>562,-8</position>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>552</ID>
<type>AE_OR2</type>
<position>709.5,-51</position>
<input>
<ID>IN_0</ID>884 </input>
<input>
<ID>IN_1</ID>885 </input>
<output>
<ID>OUT</ID>830 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>689.5,-71.5</position>
<input>
<ID>IN_0</ID>835 </input>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>559,-13.5</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>170</ID>
<type>DD_KEYPAD_HEX</type>
<position>547,-6.5</position>
<output>
<ID>OUT_0</ID>230 </output>
<output>
<ID>OUT_1</ID>231 </output>
<output>
<ID>OUT_2</ID>232 </output>
<output>
<ID>OUT_3</ID>233 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 14</lparam></gate>
<gate>
<ID>176</ID>
<type>DD_KEYPAD_HEX</type>
<position>547,-19</position>
<output>
<ID>OUT_0</ID>214 </output>
<output>
<ID>OUT_1</ID>215 </output>
<output>
<ID>OUT_2</ID>228 </output>
<output>
<ID>OUT_3</ID>229 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>179</ID>
<type>BA_DECODER_2x4</type>
<position>726.5,-91.5</position>
<input>
<ID>IN_0</ID>762 </input>
<input>
<ID>IN_1</ID>1144 </input>
<output>
<ID>OUT_0</ID>836 </output>
<output>
<ID>OUT_1</ID>839 </output>
<output>
<ID>OUT_2</ID>840 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>AE_SMALL_INVERTER</type>
<position>598.5,-15.5</position>
<input>
<ID>IN_0</ID>1043 </input>
<output>
<ID>OUT_0</ID>862 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AE_SMALL_INVERTER</type>
<position>689.5,-64</position>
<input>
<ID>IN_0</ID>761 </input>
<output>
<ID>OUT_0</ID>833 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_LABEL</type>
<position>594,-8</position>
<gparam>LABEL_TEXT Control 7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>574</ID>
<type>AE_SMALL_INVERTER</type>
<position>644,-26.5</position>
<input>
<ID>IN_0</ID>1060 </input>
<output>
<ID>OUT_0</ID>863 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>732,-92.5</position>
<gparam>LABEL_TEXT nzp</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>576</ID>
<type>AA_LABEL</type>
<position>679,-33</position>
<gparam>LABEL_TEXT This negated line here so MDR doesn't get set to 0 when  tribus is off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>EE_VDD</type>
<position>621.5,-115.5</position>
<output>
<ID>OUT_0</ID>847 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>191</ID>
<type>EE_VDD</type>
<position>621.5,-92.5</position>
<output>
<ID>OUT_0</ID>848 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_REGISTER4</type>
<position>737.5,-92</position>
<input>
<ID>IN_0</ID>836 </input>
<input>
<ID>IN_1</ID>839 </input>
<input>
<ID>IN_2</ID>840 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>844 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>195</ID>
<type>EE_VDD</type>
<position>736.5,-84.5</position>
<output>
<ID>OUT_0</ID>844 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>197</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>596,-139</position>
<input>
<ID>ENABLE_0</ID>851 </input>
<input>
<ID>IN_0</ID>867 </input>
<input>
<ID>IN_1</ID>860 </input>
<input>
<ID>IN_2</ID>861 </input>
<input>
<ID>IN_3</ID>864 </input>
<input>
<ID>IN_4</ID>870 </input>
<input>
<ID>IN_5</ID>865 </input>
<input>
<ID>IN_6</ID>866 </input>
<input>
<ID>IN_7</ID>869 </input>
<output>
<ID>OUT_0</ID>1257 </output>
<output>
<ID>OUT_1</ID>1256 </output>
<output>
<ID>OUT_2</ID>1255 </output>
<output>
<ID>OUT_3</ID>1254 </output>
<output>
<ID>OUT_4</ID>1253 </output>
<output>
<ID>OUT_5</ID>1252 </output>
<output>
<ID>OUT_6</ID>1251 </output>
<output>
<ID>OUT_7</ID>1250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>694,-49.5</position>
<gparam>LABEL_TEXT LD</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>663</ID>
<type>AA_LABEL</type>
<position>431,-80</position>
<gparam>LABEL_TEXT turn tribus off to manually input using keypads</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>665</ID>
<type>AA_LABEL</type>
<position>433.5,-92</position>
<gparam>LABEL_TEXT Bits 0-1</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>666</ID>
<type>AA_LABEL</type>
<position>433.5,-84.5</position>
<gparam>LABEL_TEXT Bits 2-3</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>669</ID>
<type>AA_LABEL</type>
<position>431,-90.5</position>
<gparam>LABEL_TEXT Read output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>671</ID>
<type>AA_LABEL</type>
<position>431,-83</position>
<gparam>LABEL_TEXT Read output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>680</ID>
<type>AA_LABEL</type>
<position>430,-103.5</position>
<gparam>LABEL_TEXT turn tribus off to manually input using keypads</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>681</ID>
<type>AA_LABEL</type>
<position>625,-73</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>682</ID>
<type>AA_LABEL</type>
<position>430.5,-111.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>683</ID>
<type>AA_LABEL</type>
<position>434,-113</position>
<gparam>LABEL_TEXT R0-R3</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>684</ID>
<type>AA_LABEL</type>
<position>566.5,-44</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>685</ID>
<type>AA_LABEL</type>
<position>566.5,-45.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>686</ID>
<type>AE_REGISTER8</type>
<position>602,-29.5</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<input>
<ID>IN_3</ID>248 </input>
<input>
<ID>IN_4</ID>263 </input>
<input>
<ID>IN_5</ID>235 </input>
<input>
<ID>IN_6</ID>234 </input>
<input>
<ID>IN_7</ID>244 </input>
<output>
<ID>OUT_0</ID>867 </output>
<output>
<ID>OUT_1</ID>860 </output>
<output>
<ID>OUT_2</ID>861 </output>
<output>
<ID>OUT_3</ID>864 </output>
<output>
<ID>OUT_4</ID>870 </output>
<output>
<ID>OUT_5</ID>865 </output>
<output>
<ID>OUT_6</ID>866 </output>
<output>
<ID>OUT_7</ID>869 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1081 </input>
<input>
<ID>count_enable</ID>1043 </input>
<input>
<ID>count_up</ID>1043 </input>
<input>
<ID>load</ID>862 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 241</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_REGISTER8</type>
<position>499,-128.5</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1152 </output>
<output>
<ID>OUT_1</ID>1151 </output>
<output>
<ID>OUT_2</ID>199 </output>
<output>
<ID>OUT_3</ID>1149 </output>
<output>
<ID>OUT_4</ID>1148 </output>
<output>
<ID>OUT_5</ID>1147 </output>
<output>
<ID>OUT_6</ID>1146 </output>
<output>
<ID>OUT_7</ID>1231 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>766 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>688</ID>
<type>AE_REGISTER8</type>
<position>619,-29.5</position>
<input>
<ID>IN_0</ID>871 </input>
<input>
<ID>IN_1</ID>872 </input>
<input>
<ID>IN_2</ID>873 </input>
<input>
<ID>IN_3</ID>876 </input>
<input>
<ID>IN_4</ID>875 </input>
<input>
<ID>IN_5</ID>877 </input>
<input>
<ID>IN_6</ID>874 </input>
<input>
<ID>IN_7</ID>878 </input>
<output>
<ID>OUT_0</ID>1046 </output>
<output>
<ID>OUT_1</ID>1045 </output>
<output>
<ID>OUT_2</ID>1041 </output>
<output>
<ID>OUT_3</ID>1040 </output>
<output>
<ID>OUT_4</ID>1039 </output>
<output>
<ID>OUT_5</ID>1038 </output>
<output>
<ID>OUT_6</ID>1037 </output>
<output>
<ID>OUT_7</ID>1036 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>849 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 234</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_REGISTER8</type>
<position>499,-115.5</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1160 </output>
<output>
<ID>OUT_1</ID>1159 </output>
<output>
<ID>OUT_2</ID>1158 </output>
<output>
<ID>OUT_3</ID>1157 </output>
<output>
<ID>OUT_4</ID>1156 </output>
<output>
<ID>OUT_5</ID>1155 </output>
<output>
<ID>OUT_6</ID>1154 </output>
<output>
<ID>OUT_7</ID>1153 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>765 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_REGISTER8</type>
<position>657,-68</position>
<input>
<ID>IN_0</ID>1070 </input>
<input>
<ID>IN_1</ID>1071 </input>
<input>
<ID>IN_2</ID>1072 </input>
<input>
<ID>IN_3</ID>1073 </input>
<input>
<ID>IN_4</ID>1074 </input>
<input>
<ID>IN_5</ID>1069 </input>
<input>
<ID>IN_6</ID>1076 </input>
<input>
<ID>IN_7</ID>1075 </input>
<output>
<ID>OUT_0</ID>1054 </output>
<output>
<ID>OUT_1</ID>1053 </output>
<output>
<ID>OUT_2</ID>1052 </output>
<output>
<ID>OUT_3</ID>1051 </output>
<output>
<ID>OUT_4</ID>1050 </output>
<output>
<ID>OUT_5</ID>1049 </output>
<output>
<ID>OUT_6</ID>1048 </output>
<output>
<ID>OUT_7</ID>1047 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>863 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_RAM_8x8</type>
<position>634,-29</position>
<input>
<ID>ADDRESS_0</ID>1046 </input>
<input>
<ID>ADDRESS_1</ID>1045 </input>
<input>
<ID>ADDRESS_2</ID>1041 </input>
<input>
<ID>ADDRESS_3</ID>1040 </input>
<input>
<ID>ADDRESS_4</ID>1039 </input>
<input>
<ID>ADDRESS_5</ID>1038 </input>
<input>
<ID>ADDRESS_6</ID>1037 </input>
<input>
<ID>ADDRESS_7</ID>1036 </input>
<input>
<ID>DATA_IN_0</ID>1077 </input>
<input>
<ID>DATA_IN_1</ID>1062 </input>
<input>
<ID>DATA_IN_2</ID>1063 </input>
<input>
<ID>DATA_IN_3</ID>1064 </input>
<input>
<ID>DATA_IN_4</ID>1065 </input>
<input>
<ID>DATA_IN_5</ID>1066 </input>
<input>
<ID>DATA_IN_6</ID>1067 </input>
<input>
<ID>DATA_IN_7</ID>1068 </input>
<output>
<ID>DATA_OUT_0</ID>1077 </output>
<output>
<ID>DATA_OUT_1</ID>1062 </output>
<output>
<ID>DATA_OUT_2</ID>1063 </output>
<output>
<ID>DATA_OUT_3</ID>1064 </output>
<output>
<ID>DATA_OUT_4</ID>1065 </output>
<output>
<ID>DATA_OUT_5</ID>1066 </output>
<output>
<ID>DATA_OUT_6</ID>1067 </output>
<output>
<ID>DATA_OUT_7</ID>1068 </output>
<input>
<ID>ENABLE_0</ID>1232 </input>
<input>
<ID>write_enable</ID>1060 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 170</lparam>
<lparam>Address:1 187</lparam>
<lparam>Address:2 204</lparam>
<lparam>Address:3 221</lparam>
<lparam>Address:4 238</lparam>
<lparam>Address:5 255</lparam>
<lparam>Address:6 10</lparam>
<lparam>Address:7 11</lparam>
<lparam>Address:8 12</lparam>
<lparam>Address:9 13</lparam>
<lparam>Address:10 14</lparam>
<lparam>Address:11 15</lparam>
<lparam>Address:254 171</lparam>
<lparam>Address:255 220</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_REGISTER8</type>
<position>674.5,-68</position>
<input>
<ID>IN_0</ID>1054 </input>
<input>
<ID>IN_1</ID>1053 </input>
<input>
<ID>IN_2</ID>1052 </input>
<input>
<ID>IN_3</ID>1051 </input>
<input>
<ID>IN_4</ID>1050 </input>
<input>
<ID>IN_5</ID>1049 </input>
<input>
<ID>IN_6</ID>1048 </input>
<input>
<ID>IN_7</ID>1047 </input>
<output>
<ID>OUT_0</ID>845 </output>
<output>
<ID>OUT_1</ID>843 </output>
<output>
<ID>OUT_2</ID>842 </output>
<output>
<ID>OUT_3</ID>841 </output>
<output>
<ID>OUT_4</ID>882 </output>
<output>
<ID>OUT_5</ID>837 </output>
<output>
<ID>OUT_6</ID>835 </output>
<output>
<ID>OUT_7</ID>761 </output>
<input>
<ID>clear</ID>1059 </input>
<input>
<ID>clock</ID>1058 </input>
<input>
<ID>load</ID>838 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>694</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>435.5,-140</position>
<input>
<ID>ENABLE_0</ID>868 </input>
<output>
<ID>OUT_0</ID>1205 </output>
<output>
<ID>OUT_1</ID>1204 </output>
<output>
<ID>OUT_2</ID>1203 </output>
<output>
<ID>OUT_3</ID>1202 </output>
<output>
<ID>OUT_4</ID>1201 </output>
<output>
<ID>OUT_5</ID>1200 </output>
<output>
<ID>OUT_6</ID>1199 </output>
<output>
<ID>OUT_7</ID>1198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>695</ID>
<type>BB_CLOCK</type>
<position>451,-60.5</position>
<output>
<ID>CLK</ID>1185 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>696</ID>
<type>AA_TOGGLE</type>
<position>591,-11</position>
<output>
<ID>OUT_0</ID>1043 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_LABEL</type>
<position>587,-18.5</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>698</ID>
<type>AA_LABEL</type>
<position>588.5,-13</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>700</ID>
<type>AA_TOGGLE</type>
<position>601,-58</position>
<output>
<ID>OUT_0</ID>1059 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_LABEL</type>
<position>595.5,-55</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>703</ID>
<type>AA_LABEL</type>
<position>599.5,-21.5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>704</ID>
<type>AA_LABEL</type>
<position>622.5,-20</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>705</ID>
<type>AA_LABEL</type>
<position>634,-20.5</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>706</ID>
<type>AA_LABEL</type>
<position>657,-75</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>707</ID>
<type>AA_TOGGLE</type>
<position>432,-133.5</position>
<output>
<ID>OUT_0</ID>868 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>709</ID>
<type>AA_TOGGLE</type>
<position>648,-23.5</position>
<output>
<ID>OUT_0</ID>1060 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_LABEL</type>
<position>432,-132</position>
<gparam>LABEL_TEXT turn tribus off to manually input using keypads</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>711</ID>
<type>AA_LABEL</type>
<position>652.5,-18.5</position>
<gparam>LABEL_TEXT Write Enable = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>712</ID>
<type>AA_LABEL</type>
<position>652,-20.5</position>
<gparam>LABEL_TEXT Output Enable = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>713</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>647.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>1232 </input>
<input>
<ID>IN_0</ID>1077 </input>
<input>
<ID>IN_1</ID>1062 </input>
<input>
<ID>IN_2</ID>1063 </input>
<input>
<ID>IN_3</ID>1064 </input>
<input>
<ID>IN_4</ID>1065 </input>
<input>
<ID>IN_5</ID>1066 </input>
<input>
<ID>IN_6</ID>1067 </input>
<input>
<ID>IN_7</ID>1068 </input>
<output>
<ID>OUT_0</ID>1070 </output>
<output>
<ID>OUT_1</ID>1071 </output>
<output>
<ID>OUT_2</ID>1072 </output>
<output>
<ID>OUT_3</ID>1073 </output>
<output>
<ID>OUT_4</ID>1074 </output>
<output>
<ID>OUT_5</ID>1069 </output>
<output>
<ID>OUT_6</ID>1076 </output>
<output>
<ID>OUT_7</ID>1075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>714</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>625.5,-67.5</position>
<input>
<ID>ENABLE_0</ID>1060 </input>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1175 </input>
<input>
<ID>IN_2</ID>1174 </input>
<input>
<ID>IN_3</ID>753 </input>
<input>
<ID>IN_4</ID>1172 </input>
<input>
<ID>IN_5</ID>1171 </input>
<input>
<ID>IN_6</ID>1170 </input>
<input>
<ID>IN_7</ID>1169 </input>
<output>
<ID>OUT_0</ID>1077 </output>
<output>
<ID>OUT_1</ID>1062 </output>
<output>
<ID>OUT_2</ID>1063 </output>
<output>
<ID>OUT_3</ID>1064 </output>
<output>
<ID>OUT_4</ID>1065 </output>
<output>
<ID>OUT_5</ID>1066 </output>
<output>
<ID>OUT_6</ID>1067 </output>
<output>
<ID>OUT_7</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>715</ID>
<type>AA_LABEL</type>
<position>676,-75</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>716</ID>
<type>AA_LABEL</type>
<position>430.5,-144.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>718</ID>
<type>AA_AND2</type>
<position>597,-42</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>852 </input>
<output>
<ID>OUT</ID>1081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>719</ID>
<type>AA_AND2</type>
<position>582.5,-59.5</position>
<input>
<ID>IN_0</ID>1080 </input>
<input>
<ID>IN_1</ID>1185 </input>
<output>
<ID>OUT</ID>1058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_TOGGLE</type>
<position>576,-58.5</position>
<output>
<ID>OUT_0</ID>1080 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>721</ID>
<type>AA_TOGGLE</type>
<position>570,-41.5</position>
<output>
<ID>OUT_0</ID>832 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>722</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>636.5,-102.5</position>
<input>
<ID>ENABLE_0</ID>1087 </input>
<input>
<ID>IN_0</ID>1330 </input>
<input>
<ID>IN_1</ID>1323 </input>
<input>
<ID>IN_10</ID>1335 </input>
<input>
<ID>IN_11</ID>1336 </input>
<input>
<ID>IN_12</ID>1333 </input>
<input>
<ID>IN_13</ID>1331 </input>
<input>
<ID>IN_14</ID>1334 </input>
<input>
<ID>IN_15</ID>1338 </input>
<input>
<ID>IN_2</ID>1327 </input>
<input>
<ID>IN_3</ID>1326 </input>
<input>
<ID>IN_4</ID>1324 </input>
<input>
<ID>IN_5</ID>1325 </input>
<input>
<ID>IN_6</ID>1328 </input>
<input>
<ID>IN_7</ID>1329 </input>
<input>
<ID>IN_8</ID>1337 </input>
<input>
<ID>IN_9</ID>1332 </input>
<output>
<ID>OUT_0</ID>1105 </output>
<output>
<ID>OUT_1</ID>1106 </output>
<output>
<ID>OUT_10</ID>1115 </output>
<output>
<ID>OUT_11</ID>1116 </output>
<output>
<ID>OUT_12</ID>1117 </output>
<output>
<ID>OUT_13</ID>1118 </output>
<output>
<ID>OUT_14</ID>1119 </output>
<output>
<ID>OUT_15</ID>1120 </output>
<output>
<ID>OUT_2</ID>1107 </output>
<output>
<ID>OUT_3</ID>1108 </output>
<output>
<ID>OUT_4</ID>1109 </output>
<output>
<ID>OUT_5</ID>1110 </output>
<output>
<ID>OUT_6</ID>1111 </output>
<output>
<ID>OUT_7</ID>1112 </output>
<output>
<ID>OUT_8</ID>1113 </output>
<output>
<ID>OUT_9</ID>1114 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>723</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>636.5,-125.5</position>
<input>
<ID>ENABLE_0</ID>1086 </input>
<input>
<ID>IN_0</ID>1307 </input>
<input>
<ID>IN_1</ID>1309 </input>
<input>
<ID>IN_10</ID>1316 </input>
<input>
<ID>IN_11</ID>1318 </input>
<input>
<ID>IN_12</ID>1319 </input>
<input>
<ID>IN_13</ID>1321 </input>
<input>
<ID>IN_14</ID>1320 </input>
<input>
<ID>IN_15</ID>1322 </input>
<input>
<ID>IN_2</ID>1308 </input>
<input>
<ID>IN_3</ID>1310 </input>
<input>
<ID>IN_4</ID>1311 </input>
<input>
<ID>IN_5</ID>1312 </input>
<input>
<ID>IN_6</ID>1314 </input>
<input>
<ID>IN_7</ID>1313 </input>
<input>
<ID>IN_8</ID>1317 </input>
<input>
<ID>IN_9</ID>1315 </input>
<output>
<ID>OUT_0</ID>1089 </output>
<output>
<ID>OUT_1</ID>1097 </output>
<output>
<ID>OUT_10</ID>1094 </output>
<output>
<ID>OUT_11</ID>1102 </output>
<output>
<ID>OUT_12</ID>1095 </output>
<output>
<ID>OUT_13</ID>1103 </output>
<output>
<ID>OUT_14</ID>1096 </output>
<output>
<ID>OUT_15</ID>1104 </output>
<output>
<ID>OUT_2</ID>1090 </output>
<output>
<ID>OUT_3</ID>1098 </output>
<output>
<ID>OUT_4</ID>1091 </output>
<output>
<ID>OUT_5</ID>1099 </output>
<output>
<ID>OUT_6</ID>1092 </output>
<output>
<ID>OUT_7</ID>1100 </output>
<output>
<ID>OUT_8</ID>1093 </output>
<output>
<ID>OUT_9</ID>1101 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>724</ID>
<type>AA_LABEL</type>
<position>614,-89.5</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>725</ID>
<type>AE_REGISTER8</type>
<position>499,-102</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1168 </output>
<output>
<ID>OUT_1</ID>1167 </output>
<output>
<ID>OUT_2</ID>1166 </output>
<output>
<ID>OUT_3</ID>1165 </output>
<output>
<ID>OUT_4</ID>1164 </output>
<output>
<ID>OUT_5</ID>1163 </output>
<output>
<ID>OUT_6</ID>1162 </output>
<output>
<ID>OUT_7</ID>1161 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>764 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_REGISTER8</type>
<position>499,-89</position>
<input>
<ID>IN_0</ID>1205 </input>
<input>
<ID>IN_1</ID>1204 </input>
<input>
<ID>IN_2</ID>1203 </input>
<input>
<ID>IN_3</ID>1202 </input>
<input>
<ID>IN_4</ID>1201 </input>
<input>
<ID>IN_5</ID>1200 </input>
<input>
<ID>IN_6</ID>1199 </input>
<input>
<ID>IN_7</ID>1198 </input>
<output>
<ID>OUT_0</ID>1184 </output>
<output>
<ID>OUT_1</ID>1175 </output>
<output>
<ID>OUT_2</ID>1174 </output>
<output>
<ID>OUT_3</ID>753 </output>
<output>
<ID>OUT_4</ID>1172 </output>
<output>
<ID>OUT_5</ID>1171 </output>
<output>
<ID>OUT_6</ID>1170 </output>
<output>
<ID>OUT_7</ID>1169 </output>
<input>
<ID>clock</ID>1185 </input>
<input>
<ID>load</ID>763 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-78</position>
<input>
<ID>IN_0</ID>1169 </input>
<input>
<ID>IN_1</ID>1161 </input>
<input>
<ID>IN_2</ID>1153 </input>
<input>
<ID>IN_3</ID>1231 </input>
<output>
<ID>OUT</ID>1176 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>728</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-89</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1162 </input>
<input>
<ID>IN_2</ID>1154 </input>
<input>
<ID>IN_3</ID>1146 </input>
<output>
<ID>OUT</ID>1177 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>729</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-100</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1163 </input>
<input>
<ID>IN_2</ID>1155 </input>
<input>
<ID>IN_3</ID>1147 </input>
<output>
<ID>OUT</ID>1178 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>730</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-109.5</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1164 </input>
<input>
<ID>IN_2</ID>1156 </input>
<input>
<ID>IN_3</ID>1148 </input>
<output>
<ID>OUT</ID>1179 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>731</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-120.5</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>1165 </input>
<input>
<ID>IN_2</ID>1157 </input>
<input>
<ID>IN_3</ID>1149 </input>
<output>
<ID>OUT</ID>1180 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>732</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-131.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1166 </input>
<input>
<ID>IN_2</ID>1158 </input>
<input>
<ID>IN_3</ID>199 </input>
<output>
<ID>OUT</ID>1181 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>733</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-142</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1167 </input>
<input>
<ID>IN_2</ID>1159 </input>
<input>
<ID>IN_3</ID>1151 </input>
<output>
<ID>OUT</ID>1182 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>734</ID>
<type>AE_MUX_4x1</type>
<position>524.5,-153</position>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1168 </input>
<input>
<ID>IN_2</ID>1160 </input>
<input>
<ID>IN_3</ID>1152 </input>
<output>
<ID>OUT</ID>1183 </output>
<input>
<ID>SEL_0</ID>1186 </input>
<input>
<ID>SEL_1</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>735</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>563,-111.5</position>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1182 </input>
<input>
<ID>IN_2</ID>1181 </input>
<input>
<ID>IN_3</ID>1180 </input>
<input>
<ID>IN_4</ID>1179 </input>
<input>
<ID>IN_5</ID>1178 </input>
<input>
<ID>IN_6</ID>1177 </input>
<input>
<ID>IN_7</ID>1176 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>736</ID>
<type>DD_KEYPAD_HEX</type>
<position>463,-78</position>
<output>
<ID>OUT_0</ID>1186 </output>
<output>
<ID>OUT_1</ID>1187 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>738</ID>
<type>AA_LABEL</type>
<position>499,-82</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>739</ID>
<type>AA_LABEL</type>
<position>499,-95</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>740</ID>
<type>AA_LABEL</type>
<position>499,-108.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>741</ID>
<type>AA_LABEL</type>
<position>499,-121.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>742</ID>
<type>AA_LABEL</type>
<position>461.5,-71</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>743</ID>
<type>DD_KEYPAD_HEX</type>
<position>463,-100.5</position>
<output>
<ID>OUT_0</ID>1196 </output>
<output>
<ID>OUT_1</ID>1197 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>744</ID>
<type>AE_MUX_4x1</type>
<position>537,-78</position>
<input>
<ID>IN_0</ID>1169 </input>
<input>
<ID>IN_1</ID>1161 </input>
<input>
<ID>IN_2</ID>1153 </input>
<input>
<ID>IN_3</ID>1231 </input>
<output>
<ID>OUT</ID>1188 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>745</ID>
<type>AE_MUX_4x1</type>
<position>537,-89</position>
<input>
<ID>IN_0</ID>1170 </input>
<input>
<ID>IN_1</ID>1162 </input>
<input>
<ID>IN_2</ID>1154 </input>
<input>
<ID>IN_3</ID>1146 </input>
<output>
<ID>OUT</ID>1189 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>746</ID>
<type>AE_MUX_4x1</type>
<position>537,-100</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1163 </input>
<input>
<ID>IN_2</ID>1155 </input>
<input>
<ID>IN_3</ID>1147 </input>
<output>
<ID>OUT</ID>1190 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>AE_MUX_4x1</type>
<position>537,-109.5</position>
<input>
<ID>IN_0</ID>1172 </input>
<input>
<ID>IN_1</ID>1164 </input>
<input>
<ID>IN_2</ID>1156 </input>
<input>
<ID>IN_3</ID>1148 </input>
<output>
<ID>OUT</ID>1191 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>748</ID>
<type>AE_MUX_4x1</type>
<position>537,-120.5</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>1165 </input>
<input>
<ID>IN_2</ID>1157 </input>
<input>
<ID>IN_3</ID>1149 </input>
<output>
<ID>OUT</ID>1192 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>749</ID>
<type>AE_MUX_4x1</type>
<position>537,-131.5</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1166 </input>
<input>
<ID>IN_2</ID>1158 </input>
<input>
<ID>IN_3</ID>199 </input>
<output>
<ID>OUT</ID>1193 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>750</ID>
<type>AE_MUX_4x1</type>
<position>537,-142</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1167 </input>
<input>
<ID>IN_2</ID>1159 </input>
<input>
<ID>IN_3</ID>1151 </input>
<output>
<ID>OUT</ID>1194 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_MUX_4x1</type>
<position>537,-153</position>
<input>
<ID>IN_0</ID>1184 </input>
<input>
<ID>IN_1</ID>1168 </input>
<input>
<ID>IN_2</ID>1160 </input>
<input>
<ID>IN_3</ID>1152 </input>
<output>
<ID>OUT</ID>1195 </output>
<input>
<ID>SEL_0</ID>1196 </input>
<input>
<ID>SEL_1</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>752</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>563,-121.5</position>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1194 </input>
<input>
<ID>IN_2</ID>1193 </input>
<input>
<ID>IN_3</ID>1192 </input>
<input>
<ID>IN_4</ID>1191 </input>
<input>
<ID>IN_5</ID>1190 </input>
<input>
<ID>IN_6</ID>1189 </input>
<input>
<ID>IN_7</ID>1188 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>753</ID>
<type>AA_LABEL</type>
<position>461.5,-93</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>754</ID>
<type>DD_KEYPAD_HEX</type>
<position>478.5,-114.5</position>
<output>
<ID>OUT_0</ID>1201 </output>
<output>
<ID>OUT_1</ID>1200 </output>
<output>
<ID>OUT_2</ID>1199 </output>
<output>
<ID>OUT_3</ID>1198 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>755</ID>
<type>DD_KEYPAD_HEX</type>
<position>478.5,-127.5</position>
<output>
<ID>OUT_0</ID>1205 </output>
<output>
<ID>OUT_1</ID>1204 </output>
<output>
<ID>OUT_2</ID>1203 </output>
<output>
<ID>OUT_3</ID>1202 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>756</ID>
<type>AA_LABEL</type>
<position>479.5,-105.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>757</ID>
<type>BA_DECODER_2x4</type>
<position>484,-73.5</position>
<input>
<ID>ENABLE</ID>1210 </input>
<input>
<ID>IN_0</ID>768 </input>
<input>
<ID>IN_1</ID>767 </input>
<output>
<ID>OUT_0</ID>763 </output>
<output>
<ID>OUT_1</ID>764 </output>
<output>
<ID>OUT_2</ID>765 </output>
<output>
<ID>OUT_3</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>AA_TOGGLE</type>
<position>478,-72</position>
<output>
<ID>OUT_0</ID>1210 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>759</ID>
<type>AA_LABEL</type>
<position>475,-72</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>760</ID>
<type>DD_KEYPAD_HEX</type>
<position>478.5,-86</position>
<output>
<ID>OUT_0</ID>768 </output>
<output>
<ID>OUT_1</ID>767 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_LABEL</type>
<position>479.5,-79</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>762</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>581,-102.5</position>
<input>
<ID>ENABLE_0</ID>195 </input>
<input>
<ID>IN_0</ID>1183 </input>
<input>
<ID>IN_1</ID>1182 </input>
<input>
<ID>IN_2</ID>1181 </input>
<input>
<ID>IN_3</ID>1180 </input>
<input>
<ID>IN_4</ID>1179 </input>
<input>
<ID>IN_5</ID>1178 </input>
<input>
<ID>IN_6</ID>1177 </input>
<input>
<ID>IN_7</ID>1176 </input>
<output>
<ID>OUT_0</ID>1249 </output>
<output>
<ID>OUT_1</ID>1248 </output>
<output>
<ID>OUT_2</ID>1247 </output>
<output>
<ID>OUT_3</ID>1245 </output>
<output>
<ID>OUT_4</ID>1245 </output>
<output>
<ID>OUT_5</ID>1245 </output>
<output>
<ID>OUT_6</ID>1245 </output>
<output>
<ID>OUT_7</ID>1245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>763</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>581,-129.5</position>
<input>
<ID>ENABLE_0</ID>1214 </input>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1194 </input>
<input>
<ID>IN_2</ID>1193 </input>
<input>
<ID>IN_3</ID>1192 </input>
<input>
<ID>IN_4</ID>1191 </input>
<input>
<ID>IN_5</ID>1190 </input>
<input>
<ID>IN_6</ID>1189 </input>
<input>
<ID>IN_7</ID>1188 </input>
<output>
<ID>OUT_0</ID>1257 </output>
<output>
<ID>OUT_1</ID>1256 </output>
<output>
<ID>OUT_2</ID>1255 </output>
<output>
<ID>OUT_3</ID>1254 </output>
<output>
<ID>OUT_4</ID>1253 </output>
<output>
<ID>OUT_5</ID>1252 </output>
<output>
<ID>OUT_6</ID>1251 </output>
<output>
<ID>OUT_7</ID>1250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_LABEL</type>
<position>581,-107.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>766</ID>
<type>AA_LABEL</type>
<position>554.5,-106.5</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>767</ID>
<type>AA_LABEL</type>
<position>581,-134.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>768</ID>
<type>AA_LABEL</type>
<position>554.5,-116.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>769</ID>
<type>EE_VDD</type>
<position>581,-122.5</position>
<output>
<ID>OUT_0</ID>1214 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>770</ID>
<type>BA_DECODER_2x4</type>
<position>628,-86</position>
<input>
<ID>ENABLE</ID>1084 </input>
<input>
<ID>IN_0</ID>1085 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<output>
<ID>OUT_1</ID>1087 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>AA_TOGGLE</type>
<position>623,-84.5</position>
<output>
<ID>OUT_0</ID>1084 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>772</ID>
<type>AA_TOGGLE</type>
<position>618.5,-87.5</position>
<output>
<ID>OUT_0</ID>1085 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>774</ID>
<type>AA_LABEL</type>
<position>613.5,-87</position>
<gparam>LABEL_TEXT Select</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>775</ID>
<type>AE_FULLADDER_4BIT</type>
<position>654,-121.5</position>
<input>
<ID>IN_0</ID>1097 </input>
<input>
<ID>IN_1</ID>1098 </input>
<input>
<ID>IN_2</ID>1099 </input>
<input>
<ID>IN_3</ID>1100 </input>
<input>
<ID>IN_B_0</ID>1089 </input>
<input>
<ID>IN_B_1</ID>1090 </input>
<input>
<ID>IN_B_2</ID>1091 </input>
<input>
<ID>IN_B_3</ID>1092 </input>
<output>
<ID>OUT_0</ID>1121 </output>
<output>
<ID>OUT_1</ID>1122 </output>
<output>
<ID>OUT_2</ID>1123 </output>
<output>
<ID>OUT_3</ID>1124 </output>
<output>
<ID>carry_out</ID>1088 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>776</ID>
<type>AE_FULLADDER_4BIT</type>
<position>654,-137.5</position>
<input>
<ID>IN_0</ID>1101 </input>
<input>
<ID>IN_1</ID>1102 </input>
<input>
<ID>IN_2</ID>1103 </input>
<input>
<ID>IN_3</ID>1104 </input>
<input>
<ID>IN_B_0</ID>1093 </input>
<input>
<ID>IN_B_1</ID>1094 </input>
<input>
<ID>IN_B_2</ID>1095 </input>
<input>
<ID>IN_B_3</ID>1096 </input>
<output>
<ID>OUT_0</ID>1125 </output>
<output>
<ID>OUT_1</ID>1126 </output>
<output>
<ID>OUT_2</ID>1127 </output>
<output>
<ID>OUT_3</ID>1128 </output>
<input>
<ID>carry_in</ID>1088 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_LABEL</type>
<position>661.5,-114</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514.5,-143,534,-143</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<intersection>514.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>514.5,-143,514.5,-104</points>
<intersection>-143 1</intersection>
<intersection>-104 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-104,514.5,-104</points>
<connection>
<GID>725</GID>
<name>OUT_1</name></connection>
<intersection>514.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1168</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>515,-154,534,-154</points>
<connection>
<GID>734</GID>
<name>IN_1</name></connection>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<intersection>515 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>515,-154,515,-105</points>
<intersection>-154 2</intersection>
<intersection>-105 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-105,515,-105</points>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection>
<intersection>515 4</intersection></hsegment></shape></wire>
<wire>
<ID>1169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>515.5,-157.5,571.5,-157.5</points>
<intersection>515.5 5</intersection>
<intersection>571.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>571.5,-157.5,571.5,-64</points>
<intersection>-157.5 1</intersection>
<intersection>-64 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>515.5,-157.5,515.5,-81</points>
<intersection>-157.5 1</intersection>
<intersection>-85 9</intersection>
<intersection>-81 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>571.5,-64,623.5,-64</points>
<connection>
<GID>714</GID>
<name>IN_7</name></connection>
<intersection>571.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>515.5,-81,534,-81</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>515.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>503,-85,515.5,-85</points>
<connection>
<GID>726</GID>
<name>OUT_7</name></connection>
<intersection>515.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516,-158,572,-158</points>
<intersection>516 7</intersection>
<intersection>572 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>572,-158,572,-65</points>
<intersection>-158 1</intersection>
<intersection>-65 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>572,-65,623.5,-65</points>
<connection>
<GID>714</GID>
<name>IN_6</name></connection>
<intersection>572 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>516,-158,516,-86</points>
<intersection>-158 1</intersection>
<intersection>-92 11</intersection>
<intersection>-86 12</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>516,-92,534,-92</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>516 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>503,-86,516,-86</points>
<connection>
<GID>726</GID>
<name>OUT_6</name></connection>
<intersection>516 7</intersection></hsegment></shape></wire>
<wire>
<ID>1171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>516.5,-158.5,572.5,-158.5</points>
<intersection>516.5 8</intersection>
<intersection>572.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>572.5,-158.5,572.5,-66</points>
<intersection>-158.5 1</intersection>
<intersection>-66 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>572.5,-66,623.5,-66</points>
<connection>
<GID>714</GID>
<name>IN_5</name></connection>
<intersection>572.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>516.5,-158.5,516.5,-87</points>
<intersection>-158.5 1</intersection>
<intersection>-103 10</intersection>
<intersection>-87 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>516.5,-103,534,-103</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>516.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>503,-87,516.5,-87</points>
<connection>
<GID>726</GID>
<name>OUT_5</name></connection>
<intersection>516.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>517,-159,573,-159</points>
<intersection>517 13</intersection>
<intersection>573 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>573,-159,573,-67</points>
<intersection>-159 1</intersection>
<intersection>-67 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>573,-67,623.5,-67</points>
<connection>
<GID>714</GID>
<name>IN_4</name></connection>
<intersection>573 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>517,-159,517,-88</points>
<intersection>-159 1</intersection>
<intersection>-112.5 16</intersection>
<intersection>-88 17</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>517,-112.5,534,-112.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>517 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>503,-88,517,-88</points>
<connection>
<GID>726</GID>
<name>OUT_4</name></connection>
<intersection>517 13</intersection></hsegment></shape></wire>
<wire>
<ID>1174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518,-160,574,-160</points>
<intersection>518 4</intersection>
<intersection>574 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>574,-160,574,-69</points>
<intersection>-160 1</intersection>
<intersection>-69 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>518,-160,518,-90</points>
<intersection>-160 1</intersection>
<intersection>-134.5 7</intersection>
<intersection>-90 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>574,-69,623.5,-69</points>
<connection>
<GID>714</GID>
<name>IN_2</name></connection>
<intersection>574 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>518,-134.5,534,-134.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>518 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>503,-90,518,-90</points>
<connection>
<GID>726</GID>
<name>OUT_2</name></connection>
<intersection>518 4</intersection></hsegment></shape></wire>
<wire>
<ID>1175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>518.5,-160.5,574.5,-160.5</points>
<intersection>518.5 8</intersection>
<intersection>574.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>574.5,-160.5,574.5,-70</points>
<intersection>-160.5 1</intersection>
<intersection>-70 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>574.5,-70,623.5,-70</points>
<connection>
<GID>714</GID>
<name>IN_1</name></connection>
<intersection>574.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>518.5,-160.5,518.5,-91</points>
<intersection>-160.5 1</intersection>
<intersection>-145 10</intersection>
<intersection>-91 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>518.5,-145,534,-145</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>518.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>503,-91,518.5,-91</points>
<connection>
<GID>726</GID>
<name>OUT_1</name></connection>
<intersection>518.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-107.5,546,-78</points>
<intersection>-107.5 2</intersection>
<intersection>-99 3</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-78,546,-78</points>
<connection>
<GID>727</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-107.5,558,-107.5</points>
<connection>
<GID>735</GID>
<name>IN_7</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>546,-99,579,-99</points>
<connection>
<GID>762</GID>
<name>IN_7</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>1177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-108.5,546,-89</points>
<intersection>-108.5 2</intersection>
<intersection>-103.5 4</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-89,546,-89</points>
<connection>
<GID>728</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-108.5,558,-108.5</points>
<connection>
<GID>735</GID>
<name>IN_6</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>546,-103.5,579,-103.5</points>
<intersection>546 0</intersection>
<intersection>579 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>579,-103.5,579,-100</points>
<connection>
<GID>762</GID>
<name>IN_6</name></connection>
<intersection>-103.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>1178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-109.5,546,-100</points>
<intersection>-109.5 2</intersection>
<intersection>-101 3</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-100,546,-100</points>
<connection>
<GID>729</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-109.5,558,-109.5</points>
<connection>
<GID>735</GID>
<name>IN_5</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>546,-101,579,-101</points>
<connection>
<GID>762</GID>
<name>IN_5</name></connection>
<intersection>546 0</intersection></hsegment></shape></wire>
<wire>
<ID>1179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-109.5,558,-109.5</points>
<connection>
<GID>730</GID>
<name>OUT</name></connection>
<intersection>547 4</intersection>
<intersection>558 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>547,-109.5,547,-102</points>
<intersection>-109.5 1</intersection>
<intersection>-102 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>547,-102,579,-102</points>
<connection>
<GID>762</GID>
<name>IN_4</name></connection>
<intersection>547 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>558,-110.5,558,-109.5</points>
<connection>
<GID>735</GID>
<name>IN_4</name></connection>
<intersection>-109.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-120.5,546,-111.5</points>
<intersection>-120.5 1</intersection>
<intersection>-111.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-120.5,546,-120.5</points>
<connection>
<GID>731</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-111.5,558,-111.5</points>
<connection>
<GID>735</GID>
<name>IN_3</name></connection>
<intersection>546 0</intersection>
<intersection>548 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>548,-111.5,548,-103</points>
<intersection>-111.5 2</intersection>
<intersection>-103 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>548,-103,579,-103</points>
<connection>
<GID>762</GID>
<name>IN_3</name></connection>
<intersection>548 3</intersection></hsegment></shape></wire>
<wire>
<ID>1181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-131.5,546,-112.5</points>
<intersection>-131.5 1</intersection>
<intersection>-112.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-131.5,546,-131.5</points>
<connection>
<GID>732</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-112.5,558,-112.5</points>
<connection>
<GID>735</GID>
<name>IN_2</name></connection>
<intersection>546 0</intersection>
<intersection>549 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>549,-112.5,549,-104</points>
<intersection>-112.5 2</intersection>
<intersection>-104 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>549,-104,579,-104</points>
<connection>
<GID>762</GID>
<name>IN_2</name></connection>
<intersection>549 3</intersection></hsegment></shape></wire>
<wire>
<ID>1182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-142,546,-113.5</points>
<intersection>-142 1</intersection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>527.5,-142,546,-142</points>
<connection>
<GID>733</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>546,-113.5,558,-113.5</points>
<connection>
<GID>735</GID>
<name>IN_1</name></connection>
<intersection>546 0</intersection>
<intersection>550 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>550,-113.5,550,-105</points>
<intersection>-113.5 2</intersection>
<intersection>-105 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>550,-105,579,-105</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>550 3</intersection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>546,-153,546,-114.5</points>
<intersection>-153 2</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>546,-114.5,558,-114.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<intersection>546 0</intersection>
<intersection>551 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527.5,-153,546,-153</points>
<connection>
<GID>734</GID>
<name>OUT</name></connection>
<intersection>546 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>551,-114.5,551,-106</points>
<intersection>-114.5 1</intersection>
<intersection>-106 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>551,-106,579,-106</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>551 3</intersection></hsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>519,-161,575,-161</points>
<intersection>519 14</intersection>
<intersection>575 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>575,-161,575,-71</points>
<intersection>-161 1</intersection>
<intersection>-71 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>519,-161,519,-92</points>
<intersection>-161 1</intersection>
<intersection>-156 17</intersection>
<intersection>-92 18</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>575,-71,623.5,-71</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>575 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>519,-156,534,-156</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>519 14</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>503,-92,519,-92</points>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection>
<intersection>519 14</intersection></hsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-133.5,455,-60.5</points>
<connection>
<GID>695</GID>
<name>CLK</name></connection>
<intersection>-133.5 8</intersection>
<intersection>-120.5 7</intersection>
<intersection>-107 6</intersection>
<intersection>-94 5</intersection>
<intersection>-60.5 11</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>455,-94,498,-94</points>
<connection>
<GID>726</GID>
<name>clock</name></connection>
<intersection>455 0</intersection>
<intersection>497 14</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>455,-107,498,-107</points>
<connection>
<GID>725</GID>
<name>clock</name></connection>
<intersection>455 0</intersection>
<intersection>497 14</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>455,-120.5,498,-120.5</points>
<connection>
<GID>689</GID>
<name>clock</name></connection>
<intersection>455 0</intersection>
<intersection>497 14</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>455,-133.5,498,-133.5</points>
<connection>
<GID>687</GID>
<name>clock</name></connection>
<intersection>455 0</intersection>
<intersection>497 14</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>455,-60.5,579.5,-60.5</points>
<connection>
<GID>719</GID>
<name>IN_1</name></connection>
<intersection>455 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>497,-133.5,497,-94</points>
<intersection>-133.5 8</intersection>
<intersection>-120.5 7</intersection>
<intersection>-107 6</intersection>
<intersection>-94 5</intersection></vsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525.5,-148,525.5,-64</points>
<connection>
<GID>734</GID>
<name>SEL_0</name></connection>
<connection>
<GID>733</GID>
<name>SEL_0</name></connection>
<connection>
<GID>732</GID>
<name>SEL_0</name></connection>
<connection>
<GID>731</GID>
<name>SEL_0</name></connection>
<connection>
<GID>730</GID>
<name>SEL_0</name></connection>
<connection>
<GID>729</GID>
<name>SEL_0</name></connection>
<connection>
<GID>728</GID>
<name>SEL_0</name></connection>
<connection>
<GID>727</GID>
<name>SEL_0</name></connection>
<intersection>-64 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>469.5,-64,525.5,-64</points>
<intersection>469.5 22</intersection>
<intersection>525.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>469.5,-89.5,469.5,-64</points>
<intersection>-89.5 23</intersection>
<intersection>-81 27</intersection>
<intersection>-64 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>439,-89.5,469.5,-89.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>469.5 22</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>468,-81,469.5,-81</points>
<connection>
<GID>736</GID>
<name>OUT_0</name></connection>
<intersection>469.5 22</intersection></hsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,-148,524.5,-63.5</points>
<connection>
<GID>734</GID>
<name>SEL_1</name></connection>
<connection>
<GID>733</GID>
<name>SEL_1</name></connection>
<connection>
<GID>732</GID>
<name>SEL_1</name></connection>
<connection>
<GID>731</GID>
<name>SEL_1</name></connection>
<connection>
<GID>730</GID>
<name>SEL_1</name></connection>
<connection>
<GID>729</GID>
<name>SEL_1</name></connection>
<connection>
<GID>728</GID>
<name>SEL_1</name></connection>
<connection>
<GID>727</GID>
<name>SEL_1</name></connection>
<intersection>-63.5 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>469,-63.5,524.5,-63.5</points>
<intersection>469 22</intersection>
<intersection>524.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>469,-88.5,469,-63.5</points>
<intersection>-88.5 25</intersection>
<intersection>-79 23</intersection>
<intersection>-63.5 21</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>468,-79,469,-79</points>
<connection>
<GID>736</GID>
<name>OUT_1</name></connection>
<intersection>469 22</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>439,-88.5,469,-88.5</points>
<connection>
<GID>124</GID>
<name>OUT_1</name></connection>
<intersection>469 22</intersection></hsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-117.5,540.5,-78</points>
<intersection>-117.5 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-78,540.5,-78</points>
<connection>
<GID>744</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-117.5,558,-117.5</points>
<connection>
<GID>752</GID>
<name>IN_7</name></connection>
<intersection>540.5 0</intersection>
<intersection>546.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>546.5,-126,546.5,-117.5</points>
<intersection>-126 4</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>546.5,-126,579,-126</points>
<connection>
<GID>763</GID>
<name>IN_7</name></connection>
<intersection>546.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-118.5,540.5,-89</points>
<intersection>-118.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-89,540.5,-89</points>
<connection>
<GID>745</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-118.5,558,-118.5</points>
<connection>
<GID>752</GID>
<name>IN_6</name></connection>
<intersection>540.5 0</intersection>
<intersection>547 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>547,-127,547,-118.5</points>
<intersection>-127 4</intersection>
<intersection>-118.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>547,-127,579,-127</points>
<connection>
<GID>763</GID>
<name>IN_6</name></connection>
<intersection>547 3</intersection></hsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-119.5,540.5,-100</points>
<intersection>-119.5 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-100,540.5,-100</points>
<connection>
<GID>746</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-119.5,558,-119.5</points>
<connection>
<GID>752</GID>
<name>IN_5</name></connection>
<intersection>540.5 0</intersection>
<intersection>549 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>549,-128,549,-119.5</points>
<intersection>-128 4</intersection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>549,-128,579,-128</points>
<connection>
<GID>763</GID>
<name>IN_5</name></connection>
<intersection>549 3</intersection></hsegment></shape></wire>
<wire>
<ID>1191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-120.5,540.5,-109.5</points>
<intersection>-120.5 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-109.5,540.5,-109.5</points>
<connection>
<GID>747</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-120.5,558,-120.5</points>
<connection>
<GID>752</GID>
<name>IN_4</name></connection>
<intersection>540.5 0</intersection>
<intersection>550.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>550.5,-129,550.5,-120.5</points>
<intersection>-129 4</intersection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>550.5,-129,579,-129</points>
<connection>
<GID>763</GID>
<name>IN_4</name></connection>
<intersection>550.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>540.5,-121.5,558,-121.5</points>
<connection>
<GID>752</GID>
<name>IN_3</name></connection>
<intersection>540.5 2</intersection>
<intersection>552.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>540.5,-121.5,540.5,-120.5</points>
<intersection>-121.5 1</intersection>
<intersection>-120.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>540,-120.5,540.5,-120.5</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<intersection>540.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>552.5,-130,552.5,-121.5</points>
<intersection>-130 5</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>552.5,-130,579,-130</points>
<connection>
<GID>763</GID>
<name>IN_3</name></connection>
<intersection>552.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-131.5,540.5,-122.5</points>
<intersection>-131.5 1</intersection>
<intersection>-122.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-131.5,540.5,-131.5</points>
<connection>
<GID>749</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-122.5,558,-122.5</points>
<connection>
<GID>752</GID>
<name>IN_2</name></connection>
<intersection>540.5 0</intersection>
<intersection>554.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>554.5,-131,554.5,-122.5</points>
<intersection>-131 4</intersection>
<intersection>-122.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>554.5,-131,579,-131</points>
<connection>
<GID>763</GID>
<name>IN_2</name></connection>
<intersection>554.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-142,540.5,-123.5</points>
<intersection>-142 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540,-142,540.5,-142</points>
<connection>
<GID>750</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,-123.5,558,-123.5</points>
<connection>
<GID>752</GID>
<name>IN_1</name></connection>
<intersection>540.5 0</intersection>
<intersection>555.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>555.5,-132,555.5,-123.5</points>
<intersection>-132 4</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>555.5,-132,579,-132</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<intersection>555.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-153,540.5,-124.5</points>
<intersection>-153 2</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540.5,-124.5,558,-124.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection>
<intersection>556.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540,-153,540.5,-153</points>
<connection>
<GID>751</GID>
<name>OUT</name></connection>
<intersection>540.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>556.5,-133,556.5,-124.5</points>
<intersection>-133 4</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>556.5,-133,579,-133</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>556.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538,-148,538,-65</points>
<connection>
<GID>751</GID>
<name>SEL_0</name></connection>
<connection>
<GID>750</GID>
<name>SEL_0</name></connection>
<connection>
<GID>749</GID>
<name>SEL_0</name></connection>
<connection>
<GID>748</GID>
<name>SEL_0</name></connection>
<connection>
<GID>747</GID>
<name>SEL_0</name></connection>
<connection>
<GID>746</GID>
<name>SEL_0</name></connection>
<connection>
<GID>745</GID>
<name>SEL_0</name></connection>
<connection>
<GID>744</GID>
<name>SEL_0</name></connection>
<intersection>-65 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>470.5,-65,538,-65</points>
<intersection>470.5 25</intersection>
<intersection>538 0</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>470.5,-103.5,470.5,-65</points>
<intersection>-103.5 26</intersection>
<intersection>-87.5 27</intersection>
<intersection>-65 24</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>468,-103.5,470.5,-103.5</points>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection>
<intersection>470.5 25</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>439,-87.5,470.5,-87.5</points>
<connection>
<GID>124</GID>
<name>OUT_2</name></connection>
<intersection>470.5 25</intersection></hsegment></shape></wire>
<wire>
<ID>1197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,-148,537,-64.5</points>
<connection>
<GID>751</GID>
<name>SEL_1</name></connection>
<connection>
<GID>750</GID>
<name>SEL_1</name></connection>
<connection>
<GID>749</GID>
<name>SEL_1</name></connection>
<connection>
<GID>748</GID>
<name>SEL_1</name></connection>
<connection>
<GID>747</GID>
<name>SEL_1</name></connection>
<connection>
<GID>746</GID>
<name>SEL_1</name></connection>
<connection>
<GID>745</GID>
<name>SEL_1</name></connection>
<connection>
<GID>744</GID>
<name>SEL_1</name></connection>
<intersection>-64.5 30</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>470,-64.5,537,-64.5</points>
<intersection>470 31</intersection>
<intersection>537 0</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>470,-101.5,470,-64.5</points>
<intersection>-101.5 32</intersection>
<intersection>-86.5 33</intersection>
<intersection>-64.5 30</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>468,-101.5,470,-101.5</points>
<connection>
<GID>743</GID>
<name>OUT_1</name></connection>
<intersection>470 31</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>439,-86.5,470,-86.5</points>
<connection>
<GID>124</GID>
<name>OUT_3</name></connection>
<intersection>470 31</intersection></hsegment></shape></wire>
<wire>
<ID>1198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-124.5,493.5,-85</points>
<intersection>-124.5 1</intersection>
<intersection>-111.5 2</intersection>
<intersection>-98 3</intersection>
<intersection>-85 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493.5,-124.5,495,-124.5</points>
<connection>
<GID>687</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>493.5,-111.5,495,-111.5</points>
<connection>
<GID>689</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>483.5,-98,495,-98</points>
<connection>
<GID>725</GID>
<name>IN_7</name></connection>
<intersection>483.5 15</intersection>
<intersection>485.5 7</intersection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>493.5,-85,495,-85</points>
<connection>
<GID>726</GID>
<name>IN_7</name></connection>
<intersection>493.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>485.5,-136.5,485.5,-98</points>
<intersection>-136.5 8</intersection>
<intersection>-98 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>437.5,-136.5,485.5,-136.5</points>
<connection>
<GID>694</GID>
<name>OUT_7</name></connection>
<intersection>485.5 7</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>483.5,-111.5,483.5,-98</points>
<connection>
<GID>754</GID>
<name>OUT_3</name></connection>
<intersection>-98 3</intersection></vsegment></shape></wire>
<wire>
<ID>1199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,-125.5,493,-86</points>
<intersection>-125.5 4</intersection>
<intersection>-113.5 2</intersection>
<intersection>-112.5 3</intersection>
<intersection>-99 5</intersection>
<intersection>-86 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-113.5,493,-113.5</points>
<connection>
<GID>754</GID>
<name>OUT_2</name></connection>
<intersection>486 7</intersection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>493,-112.5,495,-112.5</points>
<connection>
<GID>689</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>493,-125.5,495,-125.5</points>
<connection>
<GID>687</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>493,-99,495,-99</points>
<connection>
<GID>725</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>493,-86,495,-86</points>
<connection>
<GID>726</GID>
<name>IN_6</name></connection>
<intersection>493 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>486,-137.5,486,-113.5</points>
<intersection>-137.5 8</intersection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>437.5,-137.5,486,-137.5</points>
<connection>
<GID>694</GID>
<name>OUT_6</name></connection>
<intersection>486 7</intersection></hsegment></shape></wire>
<wire>
<ID>1200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,-126.5,492.5,-87</points>
<intersection>-126.5 5</intersection>
<intersection>-115.5 2</intersection>
<intersection>-113.5 4</intersection>
<intersection>-100 3</intersection>
<intersection>-87 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-115.5,492.5,-115.5</points>
<connection>
<GID>754</GID>
<name>OUT_1</name></connection>
<intersection>486.5 7</intersection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>492.5,-100,495,-100</points>
<connection>
<GID>725</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>492.5,-113.5,495,-113.5</points>
<connection>
<GID>689</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>492.5,-126.5,495,-126.5</points>
<connection>
<GID>687</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>492.5,-87,495,-87</points>
<connection>
<GID>726</GID>
<name>IN_5</name></connection>
<intersection>492.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>486.5,-138.5,486.5,-115.5</points>
<intersection>-138.5 8</intersection>
<intersection>-115.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>437.5,-138.5,486.5,-138.5</points>
<connection>
<GID>694</GID>
<name>OUT_5</name></connection>
<intersection>486.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492,-127.5,492,-88</points>
<intersection>-127.5 5</intersection>
<intersection>-117.5 2</intersection>
<intersection>-114.5 4</intersection>
<intersection>-101 3</intersection>
<intersection>-88 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-117.5,492,-117.5</points>
<connection>
<GID>754</GID>
<name>OUT_0</name></connection>
<intersection>487 7</intersection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>492,-101,495,-101</points>
<connection>
<GID>725</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>492,-114.5,495,-114.5</points>
<connection>
<GID>689</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>492,-127.5,495,-127.5</points>
<connection>
<GID>687</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>492,-88,495,-88</points>
<connection>
<GID>726</GID>
<name>IN_4</name></connection>
<intersection>492 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>487,-139.5,487,-117.5</points>
<intersection>-139.5 8</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>437.5,-139.5,487,-139.5</points>
<connection>
<GID>694</GID>
<name>OUT_4</name></connection>
<intersection>487 7</intersection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,-128.5,491.5,-89</points>
<intersection>-128.5 4</intersection>
<intersection>-124.5 2</intersection>
<intersection>-115.5 3</intersection>
<intersection>-102 12</intersection>
<intersection>-89 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-124.5,491.5,-124.5</points>
<connection>
<GID>755</GID>
<name>OUT_3</name></connection>
<intersection>487.5 10</intersection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>491.5,-115.5,495,-115.5</points>
<connection>
<GID>689</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>491.5,-128.5,495,-128.5</points>
<connection>
<GID>687</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491.5,-89,495,-89</points>
<connection>
<GID>726</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>487.5,-140.5,487.5,-124.5</points>
<intersection>-140.5 11</intersection>
<intersection>-124.5 2</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>437.5,-140.5,487.5,-140.5</points>
<connection>
<GID>694</GID>
<name>OUT_3</name></connection>
<intersection>487.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>491.5,-102,495,-102</points>
<connection>
<GID>725</GID>
<name>IN_3</name></connection>
<intersection>491.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491,-129.5,491,-90</points>
<intersection>-129.5 1</intersection>
<intersection>-126.5 2</intersection>
<intersection>-116.5 3</intersection>
<intersection>-103 4</intersection>
<intersection>-90 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,-129.5,495,-129.5</points>
<connection>
<GID>687</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-126.5,491,-126.5</points>
<connection>
<GID>755</GID>
<name>OUT_2</name></connection>
<intersection>488 6</intersection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>491,-116.5,495,-116.5</points>
<connection>
<GID>689</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>491,-103,495,-103</points>
<connection>
<GID>725</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>491,-90,495,-90</points>
<connection>
<GID>726</GID>
<name>IN_2</name></connection>
<intersection>491 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>488,-141.5,488,-126.5</points>
<intersection>-141.5 7</intersection>
<intersection>-126.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>437.5,-141.5,488,-141.5</points>
<connection>
<GID>694</GID>
<name>OUT_2</name></connection>
<intersection>488 6</intersection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490.5,-130.5,490.5,-91</points>
<intersection>-130.5 1</intersection>
<intersection>-128.5 2</intersection>
<intersection>-117.5 3</intersection>
<intersection>-104 4</intersection>
<intersection>-91 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>490.5,-130.5,495,-130.5</points>
<connection>
<GID>687</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>483.5,-128.5,490.5,-128.5</points>
<connection>
<GID>755</GID>
<name>OUT_1</name></connection>
<intersection>488.5 6</intersection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>490.5,-117.5,495,-117.5</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490.5,-104,495,-104</points>
<connection>
<GID>725</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>490.5,-91,495,-91</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>490.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>488.5,-142.5,488.5,-128.5</points>
<intersection>-142.5 7</intersection>
<intersection>-128.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>437.5,-142.5,488.5,-142.5</points>
<connection>
<GID>694</GID>
<name>OUT_1</name></connection>
<intersection>488.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490,-131.5,490,-92</points>
<intersection>-131.5 10</intersection>
<intersection>-130.5 1</intersection>
<intersection>-118.5 3</intersection>
<intersection>-105 4</intersection>
<intersection>-92 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>483.5,-130.5,490,-130.5</points>
<connection>
<GID>755</GID>
<name>OUT_0</name></connection>
<intersection>489 6</intersection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>490,-118.5,495,-118.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>490,-105,495,-105</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>490,-92,495,-92</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>489,-143.5,489,-130.5</points>
<intersection>-143.5 7</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>437.5,-143.5,489,-143.5</points>
<connection>
<GID>694</GID>
<name>OUT_0</name></connection>
<intersection>489 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>490,-131.5,495,-131.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>490 0</intersection></hsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>480,-72,481,-72</points>
<connection>
<GID>757</GID>
<name>ENABLE</name></connection>
<connection>
<GID>758</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>581,-124.5,581,-123.5</points>
<connection>
<GID>763</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>769</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-85,437,-46</points>
<connection>
<GID>124</GID>
<name>ENABLE_0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>437,-46,712.5,-46</points>
<intersection>437 0</intersection>
<intersection>712.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>712.5,-51,712.5,-46</points>
<connection>
<GID>552</GID>
<name>OUT</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>419,-195,743.5,-195</points>
<intersection>419 3</intersection>
<intersection>743.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>743.5,-195,743.5,-57.5</points>
<intersection>-195 1</intersection>
<intersection>-57.5 4</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>419,-195,419,-105.5</points>
<intersection>-195 1</intersection>
<intersection>-105.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>712.5,-57.5,743.5,-57.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>743.5 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>419,-105.5,437,-105.5</points>
<connection>
<GID>129</GID>
<name>ENABLE_0</name></connection>
<intersection>419 3</intersection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>572,-41,594,-41</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<intersection>572 5</intersection>
<intersection>578.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>578.5,-41,578.5,-38</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>572,-41.5,572,-41</points>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>691.5,-64,691.5,-64</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,-77,680.5,-62</points>
<intersection>-77 2</intersection>
<intersection>-71.5 3</intersection>
<intersection>-66 4</intersection>
<intersection>-65 1</intersection>
<intersection>-62 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>678.5,-65,680.5,-65</points>
<connection>
<GID>692</GID>
<name>OUT_6</name></connection>
<intersection>680.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>680.5,-77,691.5,-77</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>680.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>680.5,-71.5,687.5,-71.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>680.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>680.5,-66,691.5,-66</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>680.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>680.5,-62,684,-62</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>729.5,-93,733.5,-93</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<connection>
<GID>193</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680,-66,680,-58.5</points>
<intersection>-66 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680,-58.5,691.5,-58.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>680 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>678.5,-66,680,-66</points>
<connection>
<GID>692</GID>
<name>OUT_5</name></connection>
<intersection>680 0</intersection></hsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673.5,-62,673.5,-60.5</points>
<connection>
<GID>692</GID>
<name>load</name></connection>
<connection>
<GID>832</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>729.5,-92,733.5,-92</points>
<connection>
<GID>179</GID>
<name>OUT_1</name></connection>
<connection>
<GID>193</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>729.5,-91,733.5,-91</points>
<connection>
<GID>179</GID>
<name>OUT_2</name></connection>
<connection>
<GID>193</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-112,592.5,-77.5</points>
<intersection>-112 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,-112,593.5,-112</points>
<connection>
<GID>156</GID>
<name>IN_6</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>592.5,-77.5,678.5,-77.5</points>
<intersection>592.5 0</intersection>
<intersection>678.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>678.5,-77.5,678.5,-68</points>
<connection>
<GID>692</GID>
<name>OUT_3</name></connection>
<intersection>-77.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1231</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>503.5,-75,534,-75</points>
<connection>
<GID>727</GID>
<name>IN_3</name></connection>
<connection>
<GID>744</GID>
<name>IN_3</name></connection>
<intersection>503.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>503.5,-124.5,503.5,-75</points>
<intersection>-124.5 5</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-124.5,503.5,-124.5</points>
<connection>
<GID>687</GID>
<name>OUT_7</name></connection>
<intersection>503.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591.5,-113,591.5,-77</points>
<intersection>-113 1</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591.5,-113,593.5,-113</points>
<connection>
<GID>156</GID>
<name>IN_5</name></connection>
<intersection>591.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>591.5,-77,678.5,-77</points>
<intersection>591.5 0</intersection>
<intersection>678.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>678.5,-77,678.5,-69</points>
<connection>
<GID>692</GID>
<name>OUT_2</name></connection>
<intersection>-77 2</intersection></vsegment></shape></wire>
<wire>
<ID>1232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>650,-62.5,650,-29.5</points>
<intersection>-62.5 3</intersection>
<intersection>-48.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639,-29.5,650,-29.5</points>
<connection>
<GID>691</GID>
<name>ENABLE_0</name></connection>
<intersection>650 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>647.5,-48.5,650,-48.5</points>
<connection>
<GID>826</GID>
<name>OUT_0</name></connection>
<intersection>650 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>647.5,-62.5,650,-62.5</points>
<connection>
<GID>713</GID>
<name>ENABLE_0</name></connection>
<intersection>650 0</intersection></hsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,-114,590.5,-70</points>
<intersection>-114 1</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,-114,593.5,-114</points>
<connection>
<GID>156</GID>
<name>IN_4</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>590.5,-70,678.5,-70</points>
<connection>
<GID>692</GID>
<name>OUT_1</name></connection>
<intersection>590.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>736.5,-87,736.5,-85.5</points>
<connection>
<GID>193</GID>
<name>load</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,-115,589.5,-71</points>
<intersection>-115 1</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,-115,593.5,-115</points>
<connection>
<GID>156</GID>
<name>IN_3</name></connection>
<intersection>589.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,-71,678.5,-71</points>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621.5,-116.5,621.5,-116.5</points>
<connection>
<GID>834</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621.5,-93.5,621.5,-93.5</points>
<connection>
<GID>833</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>613.5,-38,613.5,-23.5</points>
<intersection>-38 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582.5,-38,613.5,-38</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<intersection>613.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>613.5,-23.5,618,-23.5</points>
<connection>
<GID>688</GID>
<name>load</name></connection>
<intersection>613.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>528,-133.5,528,11</points>
<intersection>-133.5 4</intersection>
<intersection>-109.5 5</intersection>
<intersection>-56.5 14</intersection>
<intersection>11 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>528,-133.5,596,-133.5</points>
<intersection>528 0</intersection>
<intersection>596 12</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>528,-109.5,595.5,-109.5</points>
<connection>
<GID>156</GID>
<name>ENABLE_0</name></connection>
<intersection>528 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>528,11,607,11</points>
<intersection>528 0</intersection>
<intersection>597.5 18</intersection>
<intersection>607 13</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>596,-134,596,-133.5</points>
<connection>
<GID>197</GID>
<name>ENABLE_0</name></connection>
<intersection>-133.5 4</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>607,-0.5,607,11</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>11 8</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>528,-56.5,691,-56.5</points>
<intersection>528 0</intersection>
<intersection>691 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>691,-61,691,-55.5</points>
<intersection>-61 17</intersection>
<intersection>-56.5 14</intersection>
<intersection>-55.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>691,-55.5,691.5,-55.5</points>
<connection>
<GID>140</GID>
<name>ENABLE</name></connection>
<intersection>691 15</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>690,-61,691,-61</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>691 15</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>597.5,9,597.5,11</points>
<connection>
<GID>542</GID>
<name>ENABLE_0</name></connection>
<intersection>11 8</intersection></vsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,-43,594,-43</points>
<connection>
<GID>718</GID>
<name>IN_1</name></connection>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,-101,619.5,-101</points>
<connection>
<GID>833</GID>
<name>IN_9</name></connection>
<connection>
<GID>762</GID>
<name>OUT_5</name></connection>
<intersection>583 6</intersection>
<intersection>612 10</intersection>
<intersection>613 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>613,-124,613,-101</points>
<intersection>-124 4</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>602.5,-124,619.5,-124</points>
<connection>
<GID>834</GID>
<name>IN_9</name></connection>
<intersection>602.5 7</intersection>
<intersection>613 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>583,-102,583,-101</points>
<connection>
<GID>762</GID>
<name>OUT_4</name></connection>
<intersection>-101 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>602.5,-126,602.5,-95</points>
<intersection>-126 33</intersection>
<intersection>-124 4</intersection>
<intersection>-122 11</intersection>
<intersection>-120 18</intersection>
<intersection>-118 25</intersection>
<intersection>-112 27</intersection>
<intersection>-103 30</intersection>
<intersection>-99 26</intersection>
<intersection>-95 22</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>612,-99,619.5,-99</points>
<connection>
<GID>833</GID>
<name>IN_11</name></connection>
<intersection>612 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>612,-122,612,-99</points>
<intersection>-122 11</intersection>
<intersection>-101 1</intersection>
<intersection>-99 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>602.5,-122,619.5,-122</points>
<connection>
<GID>834</GID>
<name>IN_11</name></connection>
<intersection>602.5 7</intersection>
<intersection>612 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>611,-97,619.5,-97</points>
<connection>
<GID>833</GID>
<name>IN_13</name></connection>
<intersection>611 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>611,-120,611,-97</points>
<intersection>-120 18</intersection>
<intersection>-100 19</intersection>
<intersection>-97 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>602.5,-120,619.5,-120</points>
<connection>
<GID>834</GID>
<name>IN_13</name></connection>
<intersection>602.5 7</intersection>
<intersection>611 17</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>583,-100,611,-100</points>
<connection>
<GID>762</GID>
<name>OUT_6</name></connection>
<intersection>611 17</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>602.5,-95,619.5,-95</points>
<connection>
<GID>833</GID>
<name>IN_15</name></connection>
<intersection>602.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>602.5,-118,619.5,-118</points>
<connection>
<GID>834</GID>
<name>IN_15</name></connection>
<intersection>602.5 7</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>583,-99,602.5,-99</points>
<connection>
<GID>762</GID>
<name>OUT_7</name></connection>
<intersection>602.5 7</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>597.5,-112,602.5,-112</points>
<connection>
<GID>156</GID>
<name>OUT_6</name></connection>
<intersection>602.5 7</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>583,-103,619.5,-103</points>
<connection>
<GID>762</GID>
<name>OUT_3</name></connection>
<connection>
<GID>833</GID>
<name>IN_7</name></connection>
<intersection>602.5 7</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>602.5,-126,619.5,-126</points>
<connection>
<GID>834</GID>
<name>IN_7</name></connection>
<intersection>602.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,-105,619.5,-105</points>
<connection>
<GID>833</GID>
<name>IN_5</name></connection>
<intersection>583 7</intersection>
<intersection>601.5 9</intersection>
<intersection>615 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>615,-128,615,-105</points>
<intersection>-128 4</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>615,-128,619.5,-128</points>
<connection>
<GID>834</GID>
<name>IN_5</name></connection>
<intersection>615 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>583,-105,583,-104</points>
<connection>
<GID>762</GID>
<name>OUT_2</name></connection>
<intersection>-105 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>601.5,-113,601.5,-105</points>
<intersection>-113 10</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>597.5,-113,601.5,-113</points>
<connection>
<GID>156</GID>
<name>OUT_5</name></connection>
<intersection>601.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>1248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>586.5,-107,619.5,-107</points>
<connection>
<GID>833</GID>
<name>IN_3</name></connection>
<intersection>586.5 5</intersection>
<intersection>600 7</intersection>
<intersection>616 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>616,-130,616,-107</points>
<intersection>-130 4</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>616,-130,619.5,-130</points>
<connection>
<GID>834</GID>
<name>IN_3</name></connection>
<intersection>616 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>586.5,-107,586.5,-105</points>
<intersection>-107 1</intersection>
<intersection>-105 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-105,586.5,-105</points>
<connection>
<GID>762</GID>
<name>OUT_1</name></connection>
<intersection>586.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>600,-114,600,-107</points>
<intersection>-114 8</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>597.5,-114,600,-114</points>
<connection>
<GID>156</GID>
<name>OUT_4</name></connection>
<intersection>600 7</intersection></hsegment></shape></wire>
<wire>
<ID>1249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>586,-109,619.5,-109</points>
<connection>
<GID>833</GID>
<name>IN_1</name></connection>
<intersection>586 5</intersection>
<intersection>599 7</intersection>
<intersection>617 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>617,-132,617,-109</points>
<intersection>-132 4</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>617,-132,619.5,-132</points>
<connection>
<GID>834</GID>
<name>IN_1</name></connection>
<intersection>617 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>586,-109,586,-106</points>
<intersection>-109 1</intersection>
<intersection>-106 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-106,586,-106</points>
<connection>
<GID>762</GID>
<name>OUT_0</name></connection>
<intersection>586 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>599,-115,599,-109</points>
<intersection>-115 8</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>597.5,-115,599,-115</points>
<connection>
<GID>156</GID>
<name>OUT_3</name></connection>
<intersection>599 7</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-141.5,605.5,-12</points>
<intersection>-141.5 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-141.5,605.5,-141.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>605,-12,606,-12</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-31.5,606,-12</points>
<connection>
<GID>686</GID>
<name>OUT_1</name></connection>
<intersection>-12 2</intersection></vsegment></shape></wire>
<wire>
<ID>1250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,-119,619.5,-119</points>
<connection>
<GID>834</GID>
<name>IN_14</name></connection>
<intersection>583 5</intersection>
<intersection>609.5 6</intersection>
<intersection>610.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>610.5,-119,610.5,-96</points>
<intersection>-119 1</intersection>
<intersection>-96 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>610.5,-96,619.5,-96</points>
<connection>
<GID>833</GID>
<name>IN_14</name></connection>
<intersection>610.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>583,-126,583,-119</points>
<connection>
<GID>763</GID>
<name>OUT_7</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>609.5,-135.5,609.5,-119</points>
<intersection>-135.5 7</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>598,-135.5,609.5,-135.5</points>
<connection>
<GID>197</GID>
<name>OUT_7</name></connection>
<intersection>609.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-140.5,605.5,-11</points>
<intersection>-140.5 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-140.5,605.5,-140.5</points>
<connection>
<GID>197</GID>
<name>IN_2</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>605,-11,606,-11</points>
<connection>
<GID>546</GID>
<name>IN_2</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-30.5,606,-11</points>
<connection>
<GID>686</GID>
<name>OUT_2</name></connection>
<intersection>-11 2</intersection></vsegment></shape></wire>
<wire>
<ID>1251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583.5,-121,619.5,-121</points>
<connection>
<GID>834</GID>
<name>IN_12</name></connection>
<intersection>583.5 5</intersection>
<intersection>610.5 7</intersection>
<intersection>611.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>611.5,-121,611.5,-98</points>
<intersection>-121 1</intersection>
<intersection>-98 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>611.5,-98,619.5,-98</points>
<connection>
<GID>833</GID>
<name>IN_12</name></connection>
<intersection>611.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>583.5,-127,583.5,-121</points>
<intersection>-127 6</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-127,583.5,-127</points>
<connection>
<GID>763</GID>
<name>OUT_6</name></connection>
<intersection>583.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>610.5,-136.5,610.5,-121</points>
<intersection>-136.5 8</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>598,-136.5,610.5,-136.5</points>
<connection>
<GID>197</GID>
<name>OUT_6</name></connection>
<intersection>610.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,-23.5,596.5,-15.5</points>
<connection>
<GID>571</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>596.5,-23.5,601,-23.5</points>
<connection>
<GID>686</GID>
<name>load</name></connection>
<intersection>596.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,-123,619.5,-123</points>
<connection>
<GID>834</GID>
<name>IN_10</name></connection>
<intersection>584 5</intersection>
<intersection>611.5 7</intersection>
<intersection>612.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>612.5,-123,612.5,-100</points>
<intersection>-123 1</intersection>
<intersection>-100 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>612.5,-100,619.5,-100</points>
<connection>
<GID>833</GID>
<name>IN_10</name></connection>
<intersection>612.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>584,-128,584,-123</points>
<intersection>-128 6</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-128,584,-128</points>
<connection>
<GID>763</GID>
<name>OUT_5</name></connection>
<intersection>584 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>611.5,-137.5,611.5,-123</points>
<intersection>-137.5 8</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>598,-137.5,611.5,-137.5</points>
<connection>
<GID>197</GID>
<name>OUT_5</name></connection>
<intersection>611.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>863</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>656,-62,656,-26.5</points>
<connection>
<GID>690</GID>
<name>load</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,-26.5,656,-26.5</points>
<connection>
<GID>574</GID>
<name>OUT_0</name></connection>
<intersection>656 0</intersection></hsegment></shape></wire>
<wire>
<ID>1253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584.5,-125,619.5,-125</points>
<connection>
<GID>834</GID>
<name>IN_8</name></connection>
<intersection>584.5 5</intersection>
<intersection>612.5 7</intersection>
<intersection>613.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>613.5,-125,613.5,-102</points>
<intersection>-125 1</intersection>
<intersection>-102 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>613.5,-102,619.5,-102</points>
<connection>
<GID>833</GID>
<name>IN_8</name></connection>
<intersection>613.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>584.5,-129,584.5,-125</points>
<intersection>-129 6</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-129,584.5,-129</points>
<connection>
<GID>763</GID>
<name>OUT_4</name></connection>
<intersection>584.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>612.5,-138.5,612.5,-125</points>
<intersection>-138.5 8</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>598,-138.5,612.5,-138.5</points>
<connection>
<GID>197</GID>
<name>OUT_4</name></connection>
<intersection>612.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>864</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-139.5,605.5,-10</points>
<intersection>-139.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-139.5,605.5,-139.5</points>
<connection>
<GID>197</GID>
<name>IN_3</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>605,-10,606,-10</points>
<connection>
<GID>546</GID>
<name>IN_3</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-29.5,606,-10</points>
<connection>
<GID>686</GID>
<name>OUT_3</name></connection>
<intersection>-10 2</intersection></vsegment></shape></wire>
<wire>
<ID>1254</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-127,619.5,-127</points>
<connection>
<GID>834</GID>
<name>IN_6</name></connection>
<intersection>585 5</intersection>
<intersection>613.5 7</intersection>
<intersection>614.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>614.5,-127,614.5,-104</points>
<intersection>-127 1</intersection>
<intersection>-104 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>614.5,-104,619.5,-104</points>
<connection>
<GID>833</GID>
<name>IN_6</name></connection>
<intersection>614.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>585,-130,585,-127</points>
<intersection>-130 6</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-130,585,-130</points>
<connection>
<GID>763</GID>
<name>OUT_3</name></connection>
<intersection>585 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>613.5,-139.5,613.5,-127</points>
<intersection>-139.5 8</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>598,-139.5,613.5,-139.5</points>
<connection>
<GID>197</GID>
<name>OUT_3</name></connection>
<intersection>613.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>865</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-137.5,605.5,-8</points>
<intersection>-137.5 1</intersection>
<intersection>-8 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-137.5,605.5,-137.5</points>
<connection>
<GID>197</GID>
<name>IN_5</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>605,-8,606,-8</points>
<connection>
<GID>546</GID>
<name>IN_5</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>606,-27.5,606,-8</points>
<connection>
<GID>686</GID>
<name>OUT_5</name></connection>
<intersection>-8 7</intersection></vsegment></shape></wire>
<wire>
<ID>1255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585.5,-129,619.5,-129</points>
<connection>
<GID>834</GID>
<name>IN_4</name></connection>
<intersection>585.5 5</intersection>
<intersection>614.5 7</intersection>
<intersection>615.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>615.5,-129,615.5,-106</points>
<intersection>-129 1</intersection>
<intersection>-106 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>615.5,-106,619.5,-106</points>
<connection>
<GID>833</GID>
<name>IN_4</name></connection>
<intersection>615.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>585.5,-131,585.5,-129</points>
<intersection>-131 6</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>583,-131,585.5,-131</points>
<connection>
<GID>763</GID>
<name>OUT_2</name></connection>
<intersection>585.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>614.5,-140.5,614.5,-129</points>
<intersection>-140.5 8</intersection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>598,-140.5,614.5,-140.5</points>
<connection>
<GID>197</GID>
<name>OUT_2</name></connection>
<intersection>614.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-136.5,605.5,-7</points>
<intersection>-136.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-136.5,605.5,-136.5</points>
<connection>
<GID>197</GID>
<name>IN_6</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>605,-7,606,-7</points>
<connection>
<GID>546</GID>
<name>IN_6</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-26.5,606,-7</points>
<connection>
<GID>686</GID>
<name>OUT_6</name></connection>
<intersection>-7 2</intersection></vsegment></shape></wire>
<wire>
<ID>1256</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,-131,619.5,-131</points>
<connection>
<GID>834</GID>
<name>IN_2</name></connection>
<intersection>583 5</intersection>
<intersection>615.5 6</intersection>
<intersection>616.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>616.5,-131,616.5,-108</points>
<intersection>-131 1</intersection>
<intersection>-108 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>616.5,-108,619.5,-108</points>
<connection>
<GID>833</GID>
<name>IN_2</name></connection>
<intersection>616.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>583,-132,583,-131</points>
<connection>
<GID>763</GID>
<name>OUT_1</name></connection>
<intersection>-131 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>615.5,-141.5,615.5,-131</points>
<intersection>-141.5 7</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>598,-141.5,615.5,-141.5</points>
<connection>
<GID>197</GID>
<name>OUT_1</name></connection>
<intersection>615.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-142.5,605.5,-13</points>
<intersection>-142.5 1</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-142.5,605.5,-142.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>605,-13,606,-13</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>606,-32.5,606,-13</points>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection>
<intersection>-13 4</intersection></vsegment></shape></wire>
<wire>
<ID>868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,-135,435.5,-133.5</points>
<connection>
<GID>694</GID>
<name>ENABLE_0</name></connection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434,-133.5,435.5,-133.5</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>583,-133,619.5,-133</points>
<connection>
<GID>763</GID>
<name>OUT_0</name></connection>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<intersection>616.5 5</intersection>
<intersection>617.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>617.5,-133,617.5,-110</points>
<intersection>-133 1</intersection>
<intersection>-110 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>617.5,-110,619.5,-110</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<intersection>617.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>616.5,-142.5,616.5,-133</points>
<intersection>-142.5 6</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>598,-142.5,616.5,-142.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>616.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>869</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-135.5,605.5,-6</points>
<intersection>-135.5 1</intersection>
<intersection>-6 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-135.5,605.5,-135.5</points>
<connection>
<GID>197</GID>
<name>IN_7</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>605,-6,606,-6</points>
<connection>
<GID>546</GID>
<name>IN_7</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>606,-25.5,606,-6</points>
<connection>
<GID>686</GID>
<name>OUT_7</name></connection>
<intersection>-6 4</intersection></vsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>605.5,-138.5,605.5,-9</points>
<intersection>-138.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,-138.5,605.5,-138.5</points>
<connection>
<GID>197</GID>
<name>IN_4</name></connection>
<intersection>605.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>605,-9,606,-9</points>
<connection>
<GID>546</GID>
<name>IN_4</name></connection>
<intersection>605.5 0</intersection>
<intersection>606 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>606,-28.5,606,-9</points>
<connection>
<GID>686</GID>
<name>OUT_4</name></connection>
<intersection>-9 2</intersection></vsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>609.5,-32.5,609.5,0.5</points>
<intersection>-32.5 12</intersection>
<intersection>-13 14</intersection>
<intersection>0.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>609.5,-32.5,615,-32.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>609.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,0.5,609.5,0.5</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<intersection>609.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-13,609.5,-13</points>
<connection>
<GID>546</GID>
<name>OUT_0</name></connection>
<intersection>609.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>610,-31.5,610,1.5</points>
<intersection>-31.5 12</intersection>
<intersection>-12 14</intersection>
<intersection>1.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>610,-31.5,615,-31.5</points>
<connection>
<GID>688</GID>
<name>IN_1</name></connection>
<intersection>610 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,1.5,610,1.5</points>
<connection>
<GID>542</GID>
<name>OUT_1</name></connection>
<intersection>610 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-12,610,-12</points>
<connection>
<GID>546</GID>
<name>OUT_1</name></connection>
<intersection>610 11</intersection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>610.5,-30.5,610.5,2.5</points>
<intersection>-30.5 12</intersection>
<intersection>-11 14</intersection>
<intersection>2.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>610.5,-30.5,615,-30.5</points>
<connection>
<GID>688</GID>
<name>IN_2</name></connection>
<intersection>610.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,2.5,610.5,2.5</points>
<connection>
<GID>542</GID>
<name>OUT_2</name></connection>
<intersection>610.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-11,610.5,-11</points>
<connection>
<GID>546</GID>
<name>OUT_2</name></connection>
<intersection>610.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>612.5,-26.5,612.5,6.5</points>
<intersection>-26.5 12</intersection>
<intersection>-7 14</intersection>
<intersection>6.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>612.5,-26.5,615,-26.5</points>
<connection>
<GID>688</GID>
<name>IN_6</name></connection>
<intersection>612.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,6.5,612.5,6.5</points>
<connection>
<GID>542</GID>
<name>OUT_6</name></connection>
<intersection>612.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-7,612.5,-7</points>
<connection>
<GID>546</GID>
<name>OUT_6</name></connection>
<intersection>612.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>611.5,-28.5,611.5,4.5</points>
<intersection>-28.5 12</intersection>
<intersection>-9 14</intersection>
<intersection>4.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>611.5,-28.5,615,-28.5</points>
<connection>
<GID>688</GID>
<name>IN_4</name></connection>
<intersection>611.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,4.5,611.5,4.5</points>
<connection>
<GID>542</GID>
<name>OUT_4</name></connection>
<intersection>611.5 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-9,611.5,-9</points>
<connection>
<GID>546</GID>
<name>OUT_4</name></connection>
<intersection>611.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>611,-29.5,611,3.5</points>
<intersection>-29.5 12</intersection>
<intersection>-10 14</intersection>
<intersection>3.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>611,-29.5,615,-29.5</points>
<connection>
<GID>688</GID>
<name>IN_3</name></connection>
<intersection>611 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,3.5,611,3.5</points>
<connection>
<GID>542</GID>
<name>OUT_3</name></connection>
<intersection>611 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-10,611,-10</points>
<connection>
<GID>546</GID>
<name>OUT_3</name></connection>
<intersection>611 11</intersection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>612,-27.5,612,5.5</points>
<intersection>-27.5 12</intersection>
<intersection>-8 14</intersection>
<intersection>5.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>612,-27.5,615,-27.5</points>
<connection>
<GID>688</GID>
<name>IN_5</name></connection>
<intersection>612 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>599.5,5.5,612,5.5</points>
<connection>
<GID>542</GID>
<name>OUT_5</name></connection>
<intersection>612 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-8,612,-8</points>
<connection>
<GID>546</GID>
<name>OUT_5</name></connection>
<intersection>612 11</intersection></hsegment></shape></wire>
<wire>
<ID>878</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>613,-25.5,613,7.5</points>
<intersection>-25.5 12</intersection>
<intersection>-6 14</intersection>
<intersection>7.5 15</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>613,-25.5,615,-25.5</points>
<connection>
<GID>688</GID>
<name>IN_7</name></connection>
<intersection>613 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>609,-6,613,-6</points>
<connection>
<GID>546</GID>
<name>OUT_7</name></connection>
<intersection>613 11</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>599.5,7.5,613,7.5</points>
<connection>
<GID>542</GID>
<name>OUT_7</name></connection>
<intersection>613 11</intersection></hsegment></shape></wire>
<wire>
<ID>879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607,-4.5,607,-4.5</points>
<connection>
<GID>546</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>548</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>882</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>685,-67,685,-57.5</points>
<intersection>-67 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>685,-57.5,691.5,-57.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>685 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>678.5,-67,685,-67</points>
<connection>
<GID>692</GID>
<name>OUT_4</name></connection>
<intersection>685 0</intersection></hsegment></shape></wire>
<wire>
<ID>883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568.5,-174.5,568.5,-57.5</points>
<intersection>-174.5 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420,-174.5,568.5,-174.5</points>
<intersection>420 3</intersection>
<intersection>568.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>568.5,-57.5,702,-57.5</points>
<connection>
<GID>140</GID>
<name>OUT_1</name></connection>
<intersection>568.5 0</intersection>
<intersection>702 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>420,-174.5,420,-110</points>
<intersection>-174.5 1</intersection>
<intersection>-110 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>420,-110,435,-110</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>420 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>702,-57.5,702,-56.5</points>
<intersection>-57.5 2</intersection>
<intersection>-56.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>702,-56.5,706.5,-56.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>702 5</intersection></hsegment></shape></wire>
<wire>
<ID>884</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>568,-173.5,568,-55.5</points>
<intersection>-173.5 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421,-173.5,568,-173.5</points>
<intersection>421 3</intersection>
<intersection>568 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>568,-55.5,699,-55.5</points>
<connection>
<GID>140</GID>
<name>OUT_3</name></connection>
<intersection>568 0</intersection>
<intersection>699 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>421,-173.5,421,-89.5</points>
<intersection>-173.5 1</intersection>
<intersection>-89.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>421,-89.5,435,-89.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>421 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>699,-55.5,699,-50</points>
<intersection>-55.5 2</intersection>
<intersection>-50 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>699,-50,706.5,-50</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>699 5</intersection></hsegment></shape></wire>
<wire>
<ID>885</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699,-56.5,699,-52</points>
<intersection>-56.5 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>697.5,-56.5,699,-56.5</points>
<connection>
<GID>140</GID>
<name>OUT_2</name></connection>
<intersection>699 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>699,-52,706.5,-52</points>
<connection>
<GID>552</GID>
<name>IN_1</name></connection>
<intersection>699 0</intersection></hsegment></shape></wire>
<wire>
<ID>1307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-133,634.5,-133</points>
<connection>
<GID>834</GID>
<name>OUT_0</name></connection>
<connection>
<GID>723</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-131,634.5,-131</points>
<connection>
<GID>834</GID>
<name>OUT_2</name></connection>
<connection>
<GID>723</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-132,634.5,-132</points>
<connection>
<GID>834</GID>
<name>OUT_1</name></connection>
<connection>
<GID>723</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-130,634.5,-130</points>
<connection>
<GID>834</GID>
<name>OUT_3</name></connection>
<connection>
<GID>723</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-129,634.5,-129</points>
<connection>
<GID>834</GID>
<name>OUT_4</name></connection>
<connection>
<GID>723</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-128,634.5,-128</points>
<connection>
<GID>834</GID>
<name>OUT_5</name></connection>
<connection>
<GID>723</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1313</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-126,634.5,-126</points>
<connection>
<GID>834</GID>
<name>OUT_7</name></connection>
<connection>
<GID>723</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-127,634.5,-127</points>
<connection>
<GID>834</GID>
<name>OUT_6</name></connection>
<connection>
<GID>723</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-124,634.5,-124</points>
<connection>
<GID>834</GID>
<name>OUT_9</name></connection>
<connection>
<GID>723</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-123,634.5,-123</points>
<connection>
<GID>834</GID>
<name>OUT_10</name></connection>
<connection>
<GID>723</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1317</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-125,634.5,-125</points>
<connection>
<GID>834</GID>
<name>OUT_8</name></connection>
<connection>
<GID>723</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1318</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-122,634.5,-122</points>
<connection>
<GID>834</GID>
<name>OUT_11</name></connection>
<connection>
<GID>723</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1319</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-121,634.5,-121</points>
<connection>
<GID>834</GID>
<name>OUT_12</name></connection>
<connection>
<GID>723</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-119,634.5,-119</points>
<connection>
<GID>834</GID>
<name>OUT_14</name></connection>
<connection>
<GID>723</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-120,634.5,-120</points>
<connection>
<GID>834</GID>
<name>OUT_13</name></connection>
<connection>
<GID>723</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-118,634.5,-118</points>
<connection>
<GID>834</GID>
<name>OUT_15</name></connection>
<connection>
<GID>723</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-109,634.5,-109</points>
<connection>
<GID>833</GID>
<name>OUT_1</name></connection>
<connection>
<GID>722</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-106,634.5,-106</points>
<connection>
<GID>833</GID>
<name>OUT_4</name></connection>
<connection>
<GID>722</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-105,634.5,-105</points>
<connection>
<GID>833</GID>
<name>OUT_5</name></connection>
<connection>
<GID>722</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-107,634.5,-107</points>
<connection>
<GID>833</GID>
<name>OUT_3</name></connection>
<connection>
<GID>722</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-108,634.5,-108</points>
<connection>
<GID>833</GID>
<name>OUT_2</name></connection>
<connection>
<GID>722</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-104,634.5,-104</points>
<connection>
<GID>833</GID>
<name>OUT_6</name></connection>
<connection>
<GID>722</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-103,634.5,-103</points>
<connection>
<GID>833</GID>
<name>OUT_7</name></connection>
<connection>
<GID>722</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-110,634.5,-110</points>
<connection>
<GID>833</GID>
<name>OUT_0</name></connection>
<connection>
<GID>722</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-97,634.5,-97</points>
<connection>
<GID>833</GID>
<name>OUT_13</name></connection>
<connection>
<GID>722</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-101,634.5,-101</points>
<connection>
<GID>833</GID>
<name>OUT_9</name></connection>
<connection>
<GID>722</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-98,634.5,-98</points>
<connection>
<GID>833</GID>
<name>OUT_12</name></connection>
<connection>
<GID>722</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-96,634.5,-96</points>
<connection>
<GID>833</GID>
<name>OUT_14</name></connection>
<connection>
<GID>722</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-100,634.5,-100</points>
<connection>
<GID>833</GID>
<name>OUT_10</name></connection>
<connection>
<GID>722</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-99,634.5,-99</points>
<connection>
<GID>833</GID>
<name>OUT_11</name></connection>
<connection>
<GID>722</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1337</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-102,634.5,-102</points>
<connection>
<GID>833</GID>
<name>OUT_8</name></connection>
<connection>
<GID>722</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623.5,-95,634.5,-95</points>
<connection>
<GID>833</GID>
<name>OUT_15</name></connection>
<connection>
<GID>722</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>581,-97.5,581,-94</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>719.5,-129.5,719.5,-128</points>
<connection>
<GID>128</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>697.5,-58.5,706.5,-58.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>691.5,-71.5,691.5,-71.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-129.5,534,-129.5</points>
<connection>
<GID>687</GID>
<name>OUT_2</name></connection>
<intersection>521.5 6</intersection>
<intersection>534 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>534,-129.5,534,-128.5</points>
<connection>
<GID>749</GID>
<name>IN_3</name></connection>
<intersection>-129.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>521.5,-129.5,521.5,-128.5</points>
<connection>
<GID>732</GID>
<name>IN_3</name></connection>
<intersection>-129.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>573,-36.5,573,-24.5</points>
<intersection>-36.5 2</intersection>
<intersection>-32.5 4</intersection>
<intersection>-24.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>572,-36.5,573,-36.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>573 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-24.5,573,-24.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>573 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>573,-32.5,581,-32.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>573 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>573.5,-35.5,573.5,-23.5</points>
<intersection>-35.5 2</intersection>
<intersection>-31.5 1</intersection>
<intersection>-23.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>573.5,-31.5,581,-31.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>573.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>572,-35.5,573.5,-35.5</points>
<connection>
<GID>152</GID>
<name>OUT_1</name></connection>
<intersection>573.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-23.5,573.5,-23.5</points>
<connection>
<GID>150</GID>
<name>OUT_1</name></connection>
<intersection>573.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>574,-34.5,574,-22.5</points>
<intersection>-34.5 2</intersection>
<intersection>-30.5 1</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>574,-30.5,581,-30.5</points>
<connection>
<GID>155</GID>
<name>IN_2</name></connection>
<intersection>574 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>572,-34.5,574,-34.5</points>
<connection>
<GID>152</GID>
<name>OUT_2</name></connection>
<intersection>574 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-22.5,574,-22.5</points>
<connection>
<GID>150</GID>
<name>OUT_2</name></connection>
<intersection>574 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>574.5,-33.5,574.5,-21.5</points>
<intersection>-33.5 1</intersection>
<intersection>-29.5 2</intersection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,-33.5,574.5,-33.5</points>
<connection>
<GID>152</GID>
<name>OUT_3</name></connection>
<intersection>574.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>574.5,-29.5,581,-29.5</points>
<connection>
<GID>155</GID>
<name>IN_3</name></connection>
<intersection>574.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-21.5,574.5,-21.5</points>
<connection>
<GID>150</GID>
<name>OUT_3</name></connection>
<intersection>574.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575,-32.5,575,-20.5</points>
<intersection>-32.5 1</intersection>
<intersection>-28.5 2</intersection>
<intersection>-20.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,-32.5,575,-32.5</points>
<connection>
<GID>152</GID>
<name>OUT_4</name></connection>
<intersection>575 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>575,-28.5,581,-28.5</points>
<connection>
<GID>155</GID>
<name>IN_4</name></connection>
<intersection>575 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-20.5,575,-20.5</points>
<connection>
<GID>150</GID>
<name>OUT_4</name></connection>
<intersection>575 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575.5,-31.5,575.5,-19.5</points>
<intersection>-31.5 1</intersection>
<intersection>-27.5 2</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,-31.5,575.5,-31.5</points>
<connection>
<GID>152</GID>
<name>OUT_5</name></connection>
<intersection>575.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>575.5,-27.5,581,-27.5</points>
<connection>
<GID>155</GID>
<name>IN_5</name></connection>
<intersection>575.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-19.5,575.5,-19.5</points>
<connection>
<GID>150</GID>
<name>OUT_5</name></connection>
<intersection>575.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>576,-30.5,576,-18.5</points>
<intersection>-30.5 1</intersection>
<intersection>-26.5 2</intersection>
<intersection>-18.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,-30.5,576,-30.5</points>
<connection>
<GID>152</GID>
<name>OUT_6</name></connection>
<intersection>576 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>576,-26.5,581,-26.5</points>
<connection>
<GID>155</GID>
<name>IN_6</name></connection>
<intersection>576 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-18.5,576,-18.5</points>
<connection>
<GID>150</GID>
<name>OUT_6</name></connection>
<intersection>576 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>576.5,-29.5,576.5,-17.5</points>
<intersection>-29.5 1</intersection>
<intersection>-25.5 2</intersection>
<intersection>-17.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>572,-29.5,576.5,-29.5</points>
<connection>
<GID>152</GID>
<name>OUT_7</name></connection>
<intersection>576.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>576.5,-25.5,581,-25.5</points>
<connection>
<GID>155</GID>
<name>IN_7</name></connection>
<intersection>576.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>572,-17.5,576.5,-17.5</points>
<connection>
<GID>150</GID>
<name>OUT_7</name></connection>
<intersection>576.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>562,-10.5,562,-9</points>
<connection>
<GID>158</GID>
<name>ENABLE</name></connection>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>562,-9,577.5,-9</points>
<intersection>562 0</intersection>
<intersection>577.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>577.5,-24,577.5,-9</points>
<intersection>-24 6</intersection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>577.5,-24,583,-24</points>
<connection>
<GID>155</GID>
<name>ENABLE_0</name></connection>
<intersection>577.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>561,-13.5,562,-13.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,-28,570,-13</points>
<connection>
<GID>152</GID>
<name>ENABLE_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569,-13,570,-13</points>
<intersection>569 2</intersection>
<intersection>570 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>569,-13.5,569,-13</points>
<intersection>-13.5 3</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>568,-13.5,569,-13.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>569 2</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,-16,570,-13</points>
<connection>
<GID>150</GID>
<name>ENABLE_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569,-13,570,-13</points>
<intersection>569 2</intersection>
<intersection>570 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>569,-13,569,-12.5</points>
<intersection>-13 1</intersection>
<intersection>-12.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>568,-12.5,569,-12.5</points>
<connection>
<GID>158</GID>
<name>OUT_1</name></connection>
<intersection>569 2</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>552,-24.5,552,-22</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>552,-24.5,568,-24.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>552 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>552.5,-23.5,552.5,-20</points>
<intersection>-23.5 1</intersection>
<intersection>-20 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>552.5,-23.5,568,-23.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>552.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>552,-20,552.5,-20</points>
<connection>
<GID>176</GID>
<name>OUT_1</name></connection>
<intersection>552.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>553,-22.5,553,-18</points>
<intersection>-22.5 2</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>553,-22.5,568,-22.5</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>553 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>552,-18,553,-18</points>
<connection>
<GID>176</GID>
<name>OUT_2</name></connection>
<intersection>553 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>553.5,-21.5,553.5,-16</points>
<intersection>-21.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>553.5,-21.5,568,-21.5</points>
<connection>
<GID>150</GID>
<name>IN_3</name></connection>
<intersection>553.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>552,-16,553.5,-16</points>
<connection>
<GID>176</GID>
<name>OUT_3</name></connection>
<intersection>553.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554,-20.5,554,-9.5</points>
<intersection>-20.5 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>554,-20.5,568,-20.5</points>
<connection>
<GID>150</GID>
<name>IN_4</name></connection>
<intersection>554 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>552,-9.5,554,-9.5</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>554 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>554.5,-19.5,554.5,-7.5</points>
<intersection>-19.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>554.5,-19.5,568,-19.5</points>
<connection>
<GID>150</GID>
<name>IN_5</name></connection>
<intersection>554.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>552,-7.5,554.5,-7.5</points>
<connection>
<GID>170</GID>
<name>OUT_1</name></connection>
<intersection>554.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>555,-18.5,555,-5.5</points>
<intersection>-18.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>555,-18.5,568,-18.5</points>
<connection>
<GID>150</GID>
<name>IN_6</name></connection>
<intersection>555 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>552,-5.5,555,-5.5</points>
<connection>
<GID>170</GID>
<name>OUT_2</name></connection>
<intersection>555 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>555.5,-17.5,555.5,-3.5</points>
<intersection>-17.5 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>555.5,-17.5,568,-17.5</points>
<connection>
<GID>150</GID>
<name>IN_7</name></connection>
<intersection>555.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>552,-3.5,555.5,-3.5</points>
<connection>
<GID>170</GID>
<name>OUT_3</name></connection>
<intersection>555.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-26.5,598,-26.5</points>
<connection>
<GID>686</GID>
<name>IN_6</name></connection>
<connection>
<GID>155</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-27.5,598,-27.5</points>
<connection>
<GID>686</GID>
<name>IN_5</name></connection>
<connection>
<GID>155</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-32.5,598,-32.5</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-25.5,598,-25.5</points>
<connection>
<GID>686</GID>
<name>IN_7</name></connection>
<connection>
<GID>155</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-29.5,598,-29.5</points>
<connection>
<GID>686</GID>
<name>IN_3</name></connection>
<connection>
<GID>155</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-31.5,598,-31.5</points>
<connection>
<GID>686</GID>
<name>IN_1</name></connection>
<connection>
<GID>155</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-30.5,598,-30.5</points>
<connection>
<GID>686</GID>
<name>IN_2</name></connection>
<connection>
<GID>155</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-25.5,629,-25.5</points>
<connection>
<GID>688</GID>
<name>OUT_7</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-26.5,629,-26.5</points>
<connection>
<GID>688</GID>
<name>OUT_6</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-27.5,629,-27.5</points>
<connection>
<GID>688</GID>
<name>OUT_5</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-28.5,629,-28.5</points>
<connection>
<GID>688</GID>
<name>OUT_4</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-29.5,629,-29.5</points>
<connection>
<GID>688</GID>
<name>OUT_3</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-30.5,629,-30.5</points>
<connection>
<GID>688</GID>
<name>OUT_2</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-28.5,598,-28.5</points>
<connection>
<GID>686</GID>
<name>IN_4</name></connection>
<connection>
<GID>155</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-23.5,603,-11</points>
<connection>
<GID>686</GID>
<name>count_up</name></connection>
<intersection>-23.5 18</intersection>
<intersection>-15.5 9</intersection>
<intersection>-11 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>600.5,-15.5,603,-15.5</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>593,-11,603,-11</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>603 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>602,-23.5,603,-23.5</points>
<connection>
<GID>686</GID>
<name>count_enable</name></connection>
<intersection>603 0</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-31.5,629,-31.5</points>
<connection>
<GID>688</GID>
<name>OUT_1</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,-32.5,629,-32.5</points>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection>
<connection>
<GID>691</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-64,670.5,-64</points>
<connection>
<GID>690</GID>
<name>OUT_7</name></connection>
<connection>
<GID>692</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-65,670.5,-65</points>
<connection>
<GID>692</GID>
<name>IN_6</name></connection>
<connection>
<GID>690</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445,-162,445,-36.5</points>
<intersection>-162 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>445,-36.5,568,-36.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>445 0</intersection>
<intersection>527 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>445,-162,723,-162</points>
<intersection>445 0</intersection>
<intersection>723 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>723,-162,723,-138</points>
<intersection>-162 2</intersection>
<intersection>-138 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-138,723,-138</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>723 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>527,-36.5,527,0.5</points>
<intersection>-36.5 1</intersection>
<intersection>0.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>527,0.5,595.5,0.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>527 5</intersection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-66,670.5,-66</points>
<connection>
<GID>690</GID>
<name>OUT_5</name></connection>
<connection>
<GID>692</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-67,670.5,-67</points>
<connection>
<GID>690</GID>
<name>OUT_4</name></connection>
<connection>
<GID>692</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-68,670.5,-68</points>
<connection>
<GID>692</GID>
<name>IN_3</name></connection>
<connection>
<GID>690</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-69,670.5,-69</points>
<connection>
<GID>692</GID>
<name>IN_2</name></connection>
<connection>
<GID>690</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-70,670.5,-70</points>
<connection>
<GID>690</GID>
<name>OUT_1</name></connection>
<connection>
<GID>692</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>661,-71,670.5,-71</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<connection>
<GID>692</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1058</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,-59.5,618,-34.5</points>
<connection>
<GID>688</GID>
<name>clock</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>585.5,-59.5,668.5,-59.5</points>
<connection>
<GID>719</GID>
<name>OUT</name></connection>
<intersection>618 0</intersection>
<intersection>651 5</intersection>
<intersection>668.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>668.5,-73,668.5,-59.5</points>
<intersection>-73 9</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>651,-73,651,-59.5</points>
<intersection>-73 8</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>651,-73,656,-73</points>
<connection>
<GID>690</GID>
<name>clock</name></connection>
<intersection>651 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>668.5,-73,733,-73</points>
<connection>
<GID>692</GID>
<name>clock</name></connection>
<intersection>668.5 4</intersection>
<intersection>733 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>733,-96,733,-73</points>
<intersection>-96 13</intersection>
<intersection>-73 9</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>733,-96,736.5,-96</points>
<connection>
<GID>193</GID>
<name>clock</name></connection>
<intersection>733 12</intersection></hsegment></shape></wire>
<wire>
<ID>1059</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>603,-58,603,-34.5</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<connection>
<GID>686</GID>
<name>clear</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>603,-58,668.5,-58</points>
<intersection>603 0</intersection>
<intersection>620 3</intersection>
<intersection>651 7</intersection>
<intersection>668.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>620,-58,620,-34.5</points>
<connection>
<GID>688</GID>
<name>clear</name></connection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>668.5,-73,668.5,-58</points>
<intersection>-73 9</intersection>
<intersection>-58 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>651,-73,651,-58</points>
<intersection>-73 10</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>668.5,-73,675.5,-73</points>
<connection>
<GID>692</GID>
<name>clear</name></connection>
<intersection>668.5 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>651,-73,658,-73</points>
<connection>
<GID>690</GID>
<name>clear</name></connection>
<intersection>651 7</intersection></hsegment></shape></wire>
<wire>
<ID>1060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,-23.5,646,-23.5</points>
<connection>
<GID>709</GID>
<name>OUT_0</name></connection>
<intersection>640 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>640,-41.5,640,-23.5</points>
<intersection>-41.5 4</intersection>
<intersection>-28.5 7</intersection>
<intersection>-26.5 11</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>625.5,-41.5,647.5,-41.5</points>
<intersection>625.5 8</intersection>
<intersection>640 3</intersection>
<intersection>647.5 10</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>639,-28.5,640,-28.5</points>
<connection>
<GID>691</GID>
<name>write_enable</name></connection>
<intersection>640 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>625.5,-62.5,625.5,-41.5</points>
<connection>
<GID>714</GID>
<name>ENABLE_0</name></connection>
<intersection>-41.5 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>647.5,-42.5,647.5,-41.5</points>
<connection>
<GID>826</GID>
<name>IN_0</name></connection>
<intersection>-41.5 4</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>640,-26.5,642,-26.5</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>640 3</intersection></hsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-70,645.5,-70</points>
<connection>
<GID>714</GID>
<name>OUT_1</name></connection>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>636.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>636.5,-70,636.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_1</name></connection>
<intersection>-70 1</intersection></vsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-69,645.5,-69</points>
<connection>
<GID>714</GID>
<name>OUT_2</name></connection>
<connection>
<GID>713</GID>
<name>IN_2</name></connection>
<intersection>635.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>635.5,-69,635.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_2</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-68,645.5,-68</points>
<connection>
<GID>714</GID>
<name>OUT_3</name></connection>
<connection>
<GID>713</GID>
<name>IN_3</name></connection>
<intersection>634.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>634.5,-68,634.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_3</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-67,645.5,-67</points>
<connection>
<GID>714</GID>
<name>OUT_4</name></connection>
<connection>
<GID>713</GID>
<name>IN_4</name></connection>
<intersection>633.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>633.5,-67,633.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_4</name></connection>
<intersection>-67 1</intersection></vsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-66,645.5,-66</points>
<connection>
<GID>714</GID>
<name>OUT_5</name></connection>
<connection>
<GID>713</GID>
<name>IN_5</name></connection>
<intersection>632.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>632.5,-66,632.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_5</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-65,645.5,-65</points>
<connection>
<GID>714</GID>
<name>OUT_6</name></connection>
<connection>
<GID>713</GID>
<name>IN_6</name></connection>
<intersection>631.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>631.5,-65,631.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_6</name></connection>
<intersection>-65 1</intersection></vsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-64,645.5,-64</points>
<connection>
<GID>714</GID>
<name>OUT_7</name></connection>
<connection>
<GID>713</GID>
<name>IN_7</name></connection>
<intersection>630.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>630.5,-64,630.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_7</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-66,653,-66</points>
<connection>
<GID>713</GID>
<name>OUT_5</name></connection>
<connection>
<GID>690</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-71,653,-71</points>
<connection>
<GID>713</GID>
<name>OUT_0</name></connection>
<connection>
<GID>690</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-70,653,-70</points>
<connection>
<GID>713</GID>
<name>OUT_1</name></connection>
<connection>
<GID>690</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-69,653,-69</points>
<connection>
<GID>713</GID>
<name>OUT_2</name></connection>
<connection>
<GID>690</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-68,653,-68</points>
<connection>
<GID>713</GID>
<name>OUT_3</name></connection>
<connection>
<GID>690</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-67,653,-67</points>
<connection>
<GID>713</GID>
<name>OUT_4</name></connection>
<connection>
<GID>690</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-64,653,-64</points>
<connection>
<GID>713</GID>
<name>OUT_7</name></connection>
<connection>
<GID>690</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>649.5,-65,653,-65</points>
<connection>
<GID>713</GID>
<name>OUT_6</name></connection>
<connection>
<GID>690</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>627.5,-71,645.5,-71</points>
<connection>
<GID>714</GID>
<name>OUT_0</name></connection>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>637.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>637.5,-71,637.5,-36</points>
<connection>
<GID>691</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>691</GID>
<name>DATA_IN_0</name></connection>
<intersection>-71 1</intersection></vsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578,-58.5,579.5,-58.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<connection>
<GID>720</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>601,-42,601,-34.5</points>
<connection>
<GID>686</GID>
<name>clock</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>600,-42,601,-42</points>
<connection>
<GID>718</GID>
<name>OUT</name></connection>
<intersection>601 0</intersection></hsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>625,-84.5,625,-84.5</points>
<connection>
<GID>770</GID>
<name>ENABLE</name></connection>
<connection>
<GID>771</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>620.5,-79,676.5,-79</points>
<intersection>620.5 8</intersection>
<intersection>676.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>676.5,-130.5,676.5,-79</points>
<intersection>-130.5 18</intersection>
<intersection>-125.5 19</intersection>
<intersection>-120.5 20</intersection>
<intersection>-115.5 21</intersection>
<intersection>-110.5 22</intersection>
<intersection>-105.5 23</intersection>
<intersection>-100.5 24</intersection>
<intersection>-95.5 25</intersection>
<intersection>-79 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>620.5,-87.5,620.5,-79</points>
<intersection>-87.5 10</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>620.5,-87.5,625,-87.5</points>
<connection>
<GID>772</GID>
<name>OUT_0</name></connection>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>620.5 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>676.5,-130.5,679.5,-130.5</points>
<connection>
<GID>798</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>676.5,-125.5,679.5,-125.5</points>
<connection>
<GID>797</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>676.5,-120.5,679.5,-120.5</points>
<connection>
<GID>796</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>676.5,-115.5,679.5,-115.5</points>
<connection>
<GID>795</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>676.5,-110.5,679.5,-110.5</points>
<connection>
<GID>794</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>676.5,-105.5,679.5,-105.5</points>
<connection>
<GID>793</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>676.5,-100.5,679.5,-100.5</points>
<connection>
<GID>792</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>676.5,-95.5,679.5,-95.5</points>
<connection>
<GID>791</GID>
<name>SEL_0</name></connection>
<intersection>676.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>632,-116.5,632,-87.5</points>
<intersection>-116.5 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-87.5,632,-87.5</points>
<connection>
<GID>770</GID>
<name>OUT_0</name></connection>
<intersection>632 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632,-116.5,636.5,-116.5</points>
<connection>
<GID>723</GID>
<name>ENABLE_0</name></connection>
<intersection>632 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>636.5,-93.5,636.5,-86.5</points>
<connection>
<GID>722</GID>
<name>ENABLE_0</name></connection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,-86.5,636.5,-86.5</points>
<connection>
<GID>770</GID>
<name>OUT_1</name></connection>
<intersection>636.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>653,-129.5,653,-129.5</points>
<connection>
<GID>775</GID>
<name>carry_out</name></connection>
<connection>
<GID>776</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,-133,640,-116.5</points>
<intersection>-133 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,-116.5,650,-116.5</points>
<connection>
<GID>775</GID>
<name>IN_B_0</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-133,640,-133</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640.5,-131,640.5,-117.5</points>
<intersection>-131 2</intersection>
<intersection>-117.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640.5,-117.5,650,-117.5</points>
<connection>
<GID>775</GID>
<name>IN_B_1</name></connection>
<intersection>640.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-131,640.5,-131</points>
<connection>
<GID>723</GID>
<name>OUT_2</name></connection>
<intersection>640.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641,-129,641,-118.5</points>
<intersection>-129 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641,-118.5,650,-118.5</points>
<connection>
<GID>775</GID>
<name>IN_B_2</name></connection>
<intersection>641 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-129,641,-129</points>
<connection>
<GID>723</GID>
<name>OUT_4</name></connection>
<intersection>641 0</intersection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>641.5,-127,641.5,-119.5</points>
<intersection>-127 2</intersection>
<intersection>-119.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>641.5,-119.5,650,-119.5</points>
<connection>
<GID>775</GID>
<name>IN_B_3</name></connection>
<intersection>641.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-127,641.5,-127</points>
<connection>
<GID>723</GID>
<name>OUT_6</name></connection>
<intersection>641.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643.5,-132.5,643.5,-125</points>
<intersection>-132.5 1</intersection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643.5,-132.5,650,-132.5</points>
<connection>
<GID>776</GID>
<name>IN_B_0</name></connection>
<intersection>643.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-125,643.5,-125</points>
<connection>
<GID>723</GID>
<name>OUT_8</name></connection>
<intersection>643.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643,-133.5,643,-123</points>
<intersection>-133.5 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>643,-133.5,650,-133.5</points>
<connection>
<GID>776</GID>
<name>IN_B_1</name></connection>
<intersection>643 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-123,643,-123</points>
<connection>
<GID>723</GID>
<name>OUT_10</name></connection>
<intersection>643 0</intersection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642.5,-134.5,642.5,-121</points>
<intersection>-134.5 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642.5,-134.5,650,-134.5</points>
<connection>
<GID>776</GID>
<name>IN_B_2</name></connection>
<intersection>642.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-121,642.5,-121</points>
<connection>
<GID>723</GID>
<name>OUT_12</name></connection>
<intersection>642.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642,-135.5,642,-119</points>
<intersection>-135.5 1</intersection>
<intersection>-119 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642,-135.5,650,-135.5</points>
<connection>
<GID>776</GID>
<name>IN_B_3</name></connection>
<intersection>642 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-119,642,-119</points>
<connection>
<GID>723</GID>
<name>OUT_14</name></connection>
<intersection>642 0</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-132,644,-123.5</points>
<intersection>-132 2</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-123.5,650,-123.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-132,644,-132</points>
<connection>
<GID>723</GID>
<name>OUT_1</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-130,644,-124.5</points>
<intersection>-130 2</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-124.5,650,-124.5</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-130,644,-130</points>
<connection>
<GID>723</GID>
<name>OUT_3</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-128,644,-125.5</points>
<intersection>-128 2</intersection>
<intersection>-125.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-125.5,650,-125.5</points>
<connection>
<GID>775</GID>
<name>IN_2</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-128,644,-128</points>
<connection>
<GID>723</GID>
<name>OUT_5</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644,-126.5,644,-126</points>
<intersection>-126.5 1</intersection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644,-126.5,650,-126.5</points>
<connection>
<GID>775</GID>
<name>IN_3</name></connection>
<intersection>644 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-126,644,-126</points>
<connection>
<GID>723</GID>
<name>OUT_7</name></connection>
<intersection>644 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646,-139.5,646,-124</points>
<intersection>-139.5 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,-139.5,650,-139.5</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>646 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-124,646,-124</points>
<connection>
<GID>723</GID>
<name>OUT_9</name></connection>
<intersection>646 0</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645.5,-140.5,645.5,-122</points>
<intersection>-140.5 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645.5,-140.5,650,-140.5</points>
<connection>
<GID>776</GID>
<name>IN_1</name></connection>
<intersection>645.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-122,645.5,-122</points>
<connection>
<GID>723</GID>
<name>OUT_11</name></connection>
<intersection>645.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>645,-141.5,645,-120</points>
<intersection>-141.5 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>645,-141.5,650,-141.5</points>
<connection>
<GID>776</GID>
<name>IN_2</name></connection>
<intersection>645 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-120,645,-120</points>
<connection>
<GID>723</GID>
<name>OUT_13</name></connection>
<intersection>645 0</intersection></hsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>644.5,-142.5,644.5,-118</points>
<intersection>-142.5 1</intersection>
<intersection>-118 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>644.5,-142.5,650,-142.5</points>
<connection>
<GID>776</GID>
<name>IN_3</name></connection>
<intersection>644.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-118,644.5,-118</points>
<connection>
<GID>723</GID>
<name>OUT_15</name></connection>
<intersection>644.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-112,639.5,-110</points>
<intersection>-112 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-112,646.5,-112</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-110,639.5,-110</points>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638.5,-110,646.5,-110</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>638.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>638.5,-110,638.5,-109</points>
<connection>
<GID>722</GID>
<name>OUT_1</name></connection>
<intersection>-110 1</intersection></vsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>642,-108.5,642,-108</points>
<intersection>-108.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>642,-108.5,651.5,-108.5</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>642 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-108,642,-108</points>
<connection>
<GID>722</GID>
<name>OUT_2</name></connection>
<intersection>642 0</intersection></hsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638.5,-106.5,651.5,-106.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>638.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>638.5,-107,638.5,-106.5</points>
<connection>
<GID>722</GID>
<name>OUT_3</name></connection>
<intersection>-106.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638.5,-106,646.5,-106</points>
<connection>
<GID>722</GID>
<name>OUT_4</name></connection>
<intersection>646.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>646.5,-106,646.5,-105</points>
<connection>
<GID>785</GID>
<name>IN_1</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-105,639.5,-103</points>
<intersection>-105 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-103,646.5,-103</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-105,639.5,-105</points>
<connection>
<GID>722</GID>
<name>OUT_5</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640.5,-104,640.5,-101.5</points>
<intersection>-104 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640.5,-101.5,651.5,-101.5</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>640.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-104,640.5,-104</points>
<connection>
<GID>722</GID>
<name>OUT_6</name></connection>
<intersection>640.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,-103,640,-99.5</points>
<intersection>-103 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,-99.5,651.5,-99.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-103,640,-103</points>
<connection>
<GID>722</GID>
<name>OUT_7</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-102,639.5,-98</points>
<intersection>-102 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-98,646.5,-98</points>
<connection>
<GID>787</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-102,639.5,-102</points>
<connection>
<GID>722</GID>
<name>OUT_8</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-101,639.5,-96</points>
<intersection>-101 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-96,646.5,-96</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-101,639.5,-101</points>
<connection>
<GID>722</GID>
<name>OUT_9</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,-100,640,-94.5</points>
<intersection>-100 2</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,-94.5,651.5,-94.5</points>
<connection>
<GID>788</GID>
<name>IN_1</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-100,640,-100</points>
<connection>
<GID>722</GID>
<name>OUT_10</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,-99,640,-92.5</points>
<intersection>-99 2</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,-92.5,651.5,-92.5</points>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-99,640,-99</points>
<connection>
<GID>722</GID>
<name>OUT_11</name></connection>
<intersection>640 0</intersection></hsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-98,639.5,-91</points>
<intersection>-98 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-91,646.5,-91</points>
<connection>
<GID>789</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-98,639.5,-98</points>
<connection>
<GID>722</GID>
<name>OUT_12</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,-97,639.5,-89</points>
<intersection>-97 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639.5,-89,646.5,-89</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-97,639.5,-97</points>
<connection>
<GID>722</GID>
<name>OUT_13</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639,-96,639,-87.5</points>
<intersection>-96 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>639,-87.5,651.5,-87.5</points>
<connection>
<GID>790</GID>
<name>IN_1</name></connection>
<intersection>639 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638.5,-96,639,-96</points>
<connection>
<GID>722</GID>
<name>OUT_14</name></connection>
<intersection>639 0</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638.5,-95,638.5,-85.5</points>
<connection>
<GID>722</GID>
<name>OUT_15</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638.5,-85.5,651.5,-85.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>638.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-134,667.5,-120</points>
<intersection>-134 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-134,677.5,-134</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-120,667.5,-120</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-129,667.5,-121</points>
<intersection>-129 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-129,677.5,-129</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-121,667.5,-121</points>
<connection>
<GID>775</GID>
<name>OUT_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-124,667.5,-122</points>
<intersection>-124 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-124,677.5,-124</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-122,667.5,-122</points>
<connection>
<GID>775</GID>
<name>OUT_2</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-123,667.5,-119</points>
<intersection>-123 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-119,677.5,-119</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-123,667.5,-123</points>
<connection>
<GID>775</GID>
<name>OUT_3</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-136,667.5,-114</points>
<intersection>-136 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-114,677.5,-114</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-136,667.5,-136</points>
<connection>
<GID>776</GID>
<name>OUT_0</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-137,667.5,-109</points>
<intersection>-137 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-109,677.5,-109</points>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-137,667.5,-137</points>
<connection>
<GID>776</GID>
<name>OUT_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-138,667.5,-104</points>
<intersection>-138 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-104,677.5,-104</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-138,667.5,-138</points>
<connection>
<GID>776</GID>
<name>OUT_2</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-139,667.5,-99</points>
<intersection>-139 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>667.5,-99,677.5,-99</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>658,-139,667.5,-139</points>
<connection>
<GID>776</GID>
<name>OUT_3</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,-132,665,-111</points>
<intersection>-132 1</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>665,-132,677.5,-132</points>
<connection>
<GID>798</GID>
<name>IN_1</name></connection>
<intersection>665 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>652.5,-111,665,-111</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<intersection>665 0</intersection></hsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-127,667.5,-107.5</points>
<intersection>-127 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>657.5,-107.5,667.5,-107.5</points>
<connection>
<GID>784</GID>
<name>OUT</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>667.5,-127,677.5,-127</points>
<connection>
<GID>797</GID>
<name>IN_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,-122,665,-104</points>
<intersection>-122 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>652.5,-104,665,-104</points>
<connection>
<GID>785</GID>
<name>OUT</name></connection>
<intersection>665 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>665,-122,677.5,-122</points>
<connection>
<GID>796</GID>
<name>IN_1</name></connection>
<intersection>665 0</intersection></hsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-117,667.5,-100.5</points>
<intersection>-117 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>657.5,-100.5,667.5,-100.5</points>
<connection>
<GID>786</GID>
<name>OUT</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>667.5,-117,677.5,-117</points>
<connection>
<GID>795</GID>
<name>IN_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,-112,665,-97</points>
<intersection>-112 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>652.5,-97,665,-97</points>
<connection>
<GID>787</GID>
<name>OUT</name></connection>
<intersection>665 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>665,-112,677.5,-112</points>
<connection>
<GID>794</GID>
<name>IN_1</name></connection>
<intersection>665 0</intersection></hsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-107,667.5,-93.5</points>
<intersection>-107 2</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>657.5,-93.5,667.5,-93.5</points>
<connection>
<GID>788</GID>
<name>OUT</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>667.5,-107,677.5,-107</points>
<connection>
<GID>793</GID>
<name>IN_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,-102,665,-90</points>
<intersection>-102 2</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>652.5,-90,665,-90</points>
<connection>
<GID>789</GID>
<name>OUT</name></connection>
<intersection>665 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>665,-102,677.5,-102</points>
<connection>
<GID>792</GID>
<name>IN_1</name></connection>
<intersection>665 0</intersection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,-97,667.5,-86.5</points>
<intersection>-97 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>657.5,-86.5,667.5,-86.5</points>
<connection>
<GID>790</GID>
<name>OUT</name></connection>
<intersection>667.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>667.5,-97,677.5,-97</points>
<connection>
<GID>791</GID>
<name>IN_1</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-133,689,-119</points>
<intersection>-133 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-119,720,-119</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>689 0</intersection>
<intersection>690 7</intersection>
<intersection>712 11</intersection>
<intersection>717.5 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-133,689,-133</points>
<connection>
<GID>798</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>690,-123.5,690,-119</points>
<intersection>-123.5 8</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>690,-123.5,711,-123.5</points>
<intersection>690 7</intersection>
<intersection>711 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>711,-124,711,-123.5</points>
<connection>
<GID>809</GID>
<name>N_in2</name></connection>
<intersection>-123.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>717.5,-138,717.5,-119</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>712,-119,712,-99</points>
<intersection>-119 1</intersection>
<intersection>-99 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>712,-99,715,-99</points>
<connection>
<GID>149</GID>
<name>IN_4</name></connection>
<intersection>712 11</intersection></hsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-128,689,-118</points>
<intersection>-128 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-118,720,-118</points>
<connection>
<GID>799</GID>
<name>IN_1</name></connection>
<intersection>689 0</intersection>
<intersection>690.5 7</intersection>
<intersection>711 13</intersection>
<intersection>717 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-128,689,-128</points>
<connection>
<GID>797</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>690.5,-123,690.5,-118</points>
<intersection>-123 8</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>690.5,-123,708.5,-123</points>
<intersection>690.5 7</intersection>
<intersection>708.5 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>717,-137,717,-118</points>
<intersection>-137 11</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>717,-137,717.5,-137</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>717 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>708.5,-124,708.5,-123</points>
<connection>
<GID>808</GID>
<name>N_in2</name></connection>
<intersection>-123 8</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>711,-118,711,-98</points>
<intersection>-118 1</intersection>
<intersection>-98 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>711,-98,715,-98</points>
<connection>
<GID>149</GID>
<name>IN_5</name></connection>
<intersection>711 13</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-123,689,-117</points>
<intersection>-123 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-117,720,-117</points>
<connection>
<GID>799</GID>
<name>IN_2</name></connection>
<intersection>689 0</intersection>
<intersection>691 7</intersection>
<intersection>710 13</intersection>
<intersection>716.5 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-123,689,-123</points>
<connection>
<GID>796</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>691,-122.5,691,-117</points>
<intersection>-122.5 8</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>691,-122.5,706,-122.5</points>
<intersection>691 7</intersection>
<intersection>706 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>706,-124,706,-122.5</points>
<connection>
<GID>807</GID>
<name>N_in2</name></connection>
<intersection>-122.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>716.5,-136,716.5,-117</points>
<intersection>-136 12</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>716.5,-136,717.5,-136</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>716.5 10</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>710,-117,710,-97</points>
<intersection>-117 1</intersection>
<intersection>-97 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>710,-97,715,-97</points>
<connection>
<GID>149</GID>
<name>IN_6</name></connection>
<intersection>710 13</intersection></hsegment></shape></wire>
<wire>
<ID>1140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-118,689,-116</points>
<intersection>-118 2</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-116,720,-116</points>
<connection>
<GID>799</GID>
<name>IN_3</name></connection>
<intersection>689 0</intersection>
<intersection>691.5 8</intersection>
<intersection>709 13</intersection>
<intersection>716 11</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-118,689,-118</points>
<connection>
<GID>795</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>691.5,-122,691.5,-116</points>
<intersection>-122 9</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>691.5,-122,703.5,-122</points>
<intersection>691.5 8</intersection>
<intersection>703.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>703.5,-124,703.5,-122</points>
<connection>
<GID>806</GID>
<name>N_in2</name></connection>
<intersection>-122 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>716,-135,716,-116</points>
<intersection>-135 12</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>716,-135,717.5,-135</points>
<connection>
<GID>128</GID>
<name>IN_3</name></connection>
<intersection>716 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>709,-116,709,-96</points>
<intersection>-116 1</intersection>
<intersection>-96 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>709,-96,715,-96</points>
<connection>
<GID>149</GID>
<name>IN_7</name></connection>
<intersection>709 13</intersection></hsegment></shape></wire>
<wire>
<ID>1141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-115,689,-113</points>
<intersection>-115 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-115,720,-115</points>
<connection>
<GID>799</GID>
<name>IN_4</name></connection>
<intersection>689 0</intersection>
<intersection>692 8</intersection>
<intersection>708 13</intersection>
<intersection>715.5 11</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-113,689,-113</points>
<connection>
<GID>794</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>692,-121.5,692,-115</points>
<intersection>-121.5 9</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>692,-121.5,701,-121.5</points>
<intersection>692 8</intersection>
<intersection>701 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>701,-124,701,-121.5</points>
<connection>
<GID>805</GID>
<name>N_in2</name></connection>
<intersection>-121.5 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>715.5,-134,715.5,-115</points>
<intersection>-134 12</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>715.5,-134,717.5,-134</points>
<connection>
<GID>128</GID>
<name>IN_4</name></connection>
<intersection>715.5 11</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>708,-115,708,-95</points>
<intersection>-115 1</intersection>
<intersection>-95 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>708,-95,715,-95</points>
<connection>
<GID>149</GID>
<name>IN_3</name></connection>
<intersection>708 13</intersection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>573.5,-159.5,573.5,-68</points>
<intersection>-159.5 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>573.5,-68,623.5,-68</points>
<connection>
<GID>714</GID>
<name>IN_3</name></connection>
<intersection>573.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>517.5,-159.5,573.5,-159.5</points>
<intersection>517.5 3</intersection>
<intersection>573.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>517.5,-159.5,517.5,-89</points>
<intersection>-159.5 2</intersection>
<intersection>-123.5 6</intersection>
<intersection>-89 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-89,517.5,-89</points>
<connection>
<GID>726</GID>
<name>OUT_3</name></connection>
<intersection>517.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>517.5,-123.5,534,-123.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>517.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-114,689,-108</points>
<intersection>-114 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-114,720,-114</points>
<connection>
<GID>799</GID>
<name>IN_5</name></connection>
<intersection>689 0</intersection>
<intersection>692.5 7</intersection>
<intersection>713.5 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-108,689,-108</points>
<connection>
<GID>793</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>692.5,-121,692.5,-114</points>
<intersection>-121 8</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>692.5,-121,698.5,-121</points>
<intersection>692.5 7</intersection>
<intersection>698.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>698.5,-124,698.5,-121</points>
<connection>
<GID>804</GID>
<name>N_in2</name></connection>
<intersection>-121 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>713.5,-133,713.5,-94</points>
<intersection>-133 11</intersection>
<intersection>-114 1</intersection>
<intersection>-94 13</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>713.5,-133,717.5,-133</points>
<connection>
<GID>128</GID>
<name>IN_5</name></connection>
<intersection>713.5 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>713.5,-94,715,-94</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>713.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-113,689,-103</points>
<intersection>-113 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>689,-113,720,-113</points>
<connection>
<GID>799</GID>
<name>IN_6</name></connection>
<intersection>689 0</intersection>
<intersection>693 7</intersection>
<intersection>707 12</intersection>
<intersection>714.5 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>681.5,-103,689,-103</points>
<connection>
<GID>792</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>693,-120.5,693,-113</points>
<intersection>-120.5 8</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>693,-120.5,696,-120.5</points>
<intersection>693 7</intersection>
<intersection>696 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>696,-124,696,-120.5</points>
<connection>
<GID>803</GID>
<name>N_in2</name></connection>
<intersection>-120.5 8</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>714.5,-132,714.5,-113</points>
<intersection>-132 11</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>714.5,-132,717.5,-132</points>
<connection>
<GID>128</GID>
<name>IN_6</name></connection>
<intersection>714.5 10</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>707,-113,707,-93</points>
<intersection>-113 1</intersection>
<intersection>-93 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>707,-93,715,-93</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>707 12</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,-162.5,444.5,-35.5</points>
<intersection>-162.5 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,-35.5,568,-35.5</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>444.5 0</intersection>
<intersection>526 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444.5,-162.5,723.5,-162.5</points>
<intersection>444.5 0</intersection>
<intersection>723.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>723.5,-162.5,723.5,-137</points>
<intersection>-162.5 2</intersection>
<intersection>-137 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-137,723.5,-137</points>
<connection>
<GID>128</GID>
<name>OUT_1</name></connection>
<intersection>723.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>526,-35.5,526,1.5</points>
<intersection>-35.5 1</intersection>
<intersection>1.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>526,1.5,595.5,1.5</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>526 5</intersection></hsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,-112,689,-98</points>
<intersection>-112 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>681.5,-98,689,-98</points>
<connection>
<GID>791</GID>
<name>OUT</name></connection>
<intersection>689 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>689,-112,720,-112</points>
<connection>
<GID>799</GID>
<name>IN_7</name></connection>
<intersection>689 0</intersection>
<intersection>693.5 5</intersection>
<intersection>706 8</intersection>
<intersection>714 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>693.5,-124,693.5,-112</points>
<connection>
<GID>802</GID>
<name>N_in2</name></connection>
<intersection>-112 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>714,-131,714,-112</points>
<intersection>-131 7</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>714,-131,717.5,-131</points>
<connection>
<GID>128</GID>
<name>IN_7</name></connection>
<intersection>714 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>706,-112,706,-91</points>
<intersection>-112 2</intersection>
<intersection>-91 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>706,-91,723.5,-91</points>
<intersection>706 8</intersection>
<intersection>715 12</intersection>
<intersection>723.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>723.5,-92,723.5,-91</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>-91 9</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>715,-92,715,-91</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-91 9</intersection></vsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,-163,444,-34.5</points>
<intersection>-163 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444,-34.5,568,-34.5</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<intersection>444 0</intersection>
<intersection>525 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,-163,724,-163</points>
<intersection>444 0</intersection>
<intersection>724 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>724,-163,724,-136</points>
<intersection>-163 2</intersection>
<intersection>-136 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-136,724,-136</points>
<connection>
<GID>128</GID>
<name>OUT_2</name></connection>
<intersection>724 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>525,-34.5,525,2.5</points>
<intersection>-34.5 1</intersection>
<intersection>2.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>525,2.5,595.5,2.5</points>
<connection>
<GID>542</GID>
<name>IN_2</name></connection>
<intersection>525 5</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443.5,-163.5,443.5,-33.5</points>
<intersection>-163.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443.5,-33.5,568,-33.5</points>
<connection>
<GID>152</GID>
<name>IN_3</name></connection>
<intersection>443.5 0</intersection>
<intersection>524 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443.5,-163.5,724.5,-163.5</points>
<intersection>443.5 0</intersection>
<intersection>724.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>724.5,-163.5,724.5,-135</points>
<intersection>-163.5 2</intersection>
<intersection>-135 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-135,724.5,-135</points>
<connection>
<GID>128</GID>
<name>OUT_3</name></connection>
<intersection>724.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>524,-33.5,524,3.5</points>
<intersection>-33.5 1</intersection>
<intersection>3.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>524,3.5,595.5,3.5</points>
<connection>
<GID>542</GID>
<name>IN_3</name></connection>
<intersection>524 5</intersection></hsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-125.5,534,-125.5</points>
<connection>
<GID>687</GID>
<name>OUT_6</name></connection>
<intersection>521.5 4</intersection>
<intersection>534 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>534,-125.5,534,-86</points>
<connection>
<GID>745</GID>
<name>IN_3</name></connection>
<intersection>-125.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>521.5,-125.5,521.5,-86</points>
<connection>
<GID>728</GID>
<name>IN_3</name></connection>
<intersection>-125.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,-164,443,-32.5</points>
<intersection>-164 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443,-32.5,568,-32.5</points>
<connection>
<GID>152</GID>
<name>IN_4</name></connection>
<intersection>443 0</intersection>
<intersection>523 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443,-164,725,-164</points>
<intersection>443 0</intersection>
<intersection>725 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>725,-164,725,-134</points>
<intersection>-164 2</intersection>
<intersection>-134 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-134,725,-134</points>
<connection>
<GID>128</GID>
<name>OUT_4</name></connection>
<intersection>725 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>523,-32.5,523,4.5</points>
<intersection>-32.5 1</intersection>
<intersection>4.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>523,4.5,595.5,4.5</points>
<connection>
<GID>542</GID>
<name>IN_4</name></connection>
<intersection>523 5</intersection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>504.5,-97,534,-97</points>
<connection>
<GID>729</GID>
<name>IN_3</name></connection>
<connection>
<GID>746</GID>
<name>IN_3</name></connection>
<intersection>504.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>504.5,-126.5,504.5,-97</points>
<intersection>-126.5 5</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-126.5,504.5,-126.5</points>
<connection>
<GID>687</GID>
<name>OUT_5</name></connection>
<intersection>504.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,-164.5,442.5,-31.5</points>
<intersection>-164.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442.5,-31.5,568,-31.5</points>
<connection>
<GID>152</GID>
<name>IN_5</name></connection>
<intersection>442.5 0</intersection>
<intersection>522 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442.5,-164.5,725.5,-164.5</points>
<intersection>442.5 0</intersection>
<intersection>725.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>725.5,-164.5,725.5,-133</points>
<intersection>-164.5 2</intersection>
<intersection>-133 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-133,725.5,-133</points>
<connection>
<GID>128</GID>
<name>OUT_5</name></connection>
<intersection>725.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>522,-31.5,522,5.5</points>
<intersection>-31.5 1</intersection>
<intersection>5.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>522,5.5,595.5,5.5</points>
<connection>
<GID>542</GID>
<name>IN_5</name></connection>
<intersection>522 5</intersection></hsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>505,-106.5,534,-106.5</points>
<connection>
<GID>730</GID>
<name>IN_3</name></connection>
<connection>
<GID>747</GID>
<name>IN_3</name></connection>
<intersection>505 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>505,-127.5,505,-106.5</points>
<intersection>-127.5 6</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>503,-127.5,505,-127.5</points>
<connection>
<GID>687</GID>
<name>OUT_4</name></connection>
<intersection>505 4</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442,-165,442,-30.5</points>
<intersection>-165 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,-30.5,568,-30.5</points>
<connection>
<GID>152</GID>
<name>IN_6</name></connection>
<intersection>442 0</intersection>
<intersection>521 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442,-165,726,-165</points>
<intersection>442 0</intersection>
<intersection>726 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>726,-165,726,-132</points>
<intersection>-165 2</intersection>
<intersection>-132 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-132,726,-132</points>
<connection>
<GID>128</GID>
<name>OUT_6</name></connection>
<intersection>726 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>521,-30.5,521,6.5</points>
<intersection>-30.5 1</intersection>
<intersection>6.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>521,6.5,595.5,6.5</points>
<connection>
<GID>542</GID>
<name>IN_6</name></connection>
<intersection>521 5</intersection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>505.5,-117.5,534,-117.5</points>
<connection>
<GID>731</GID>
<name>IN_3</name></connection>
<connection>
<GID>748</GID>
<name>IN_3</name></connection>
<intersection>505.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>505.5,-128.5,505.5,-117.5</points>
<intersection>-128.5 5</intersection>
<intersection>-117.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-128.5,505.5,-128.5</points>
<connection>
<GID>687</GID>
<name>OUT_3</name></connection>
<intersection>505.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,-165.5,441.5,-29.5</points>
<intersection>-165.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,-29.5,568,-29.5</points>
<connection>
<GID>152</GID>
<name>IN_7</name></connection>
<intersection>441.5 0</intersection>
<intersection>520 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>441.5,-165.5,726.5,-165.5</points>
<intersection>441.5 0</intersection>
<intersection>726.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>726.5,-165.5,726.5,-131</points>
<intersection>-165.5 2</intersection>
<intersection>-131 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>721.5,-131,726.5,-131</points>
<connection>
<GID>128</GID>
<name>OUT_7</name></connection>
<intersection>726.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>520,-29.5,520,7.5</points>
<intersection>-29.5 1</intersection>
<intersection>7.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>520,7.5,595.5,7.5</points>
<connection>
<GID>542</GID>
<name>IN_7</name></connection>
<intersection>520 5</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>679.5,-75,679.5,-60</points>
<intersection>-75 6</intersection>
<intersection>-69.5 2</intersection>
<intersection>-64 1</intersection>
<intersection>-60 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>678.5,-64,687.5,-64</points>
<connection>
<GID>692</GID>
<name>OUT_7</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>679.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>679.5,-69.5,691.5,-69.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>679.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>679.5,-75,691.5,-75</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>679.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>679.5,-60,684,-60</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>679.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>506.5,-139,534,-139</points>
<connection>
<GID>733</GID>
<name>IN_3</name></connection>
<connection>
<GID>750</GID>
<name>IN_3</name></connection>
<intersection>506.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>506.5,-139,506.5,-130.5</points>
<intersection>-139 1</intersection>
<intersection>-130.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-130.5,506.5,-130.5</points>
<connection>
<GID>687</GID>
<name>OUT_1</name></connection>
<intersection>506.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>722.5,-95.5,722.5,-93</points>
<intersection>-95.5 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>722.5,-93,723.5,-93</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>722.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>722,-95.5,722.5,-95.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>722.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-83,497,-75</points>
<intersection>-83 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-75,497,-75</points>
<connection>
<GID>757</GID>
<name>OUT_0</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-83,498,-83</points>
<connection>
<GID>726</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1152</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>507,-150,534,-150</points>
<connection>
<GID>734</GID>
<name>IN_3</name></connection>
<connection>
<GID>751</GID>
<name>IN_3</name></connection>
<intersection>507 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>507,-150,507,-131.5</points>
<intersection>-150 2</intersection>
<intersection>-131.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-131.5,507,-131.5</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>507 4</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-96,497,-74</points>
<intersection>-96 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-74,497,-74</points>
<connection>
<GID>757</GID>
<name>OUT_1</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-96,498,-96</points>
<connection>
<GID>725</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>507.5,-77,534,-77</points>
<connection>
<GID>727</GID>
<name>IN_2</name></connection>
<connection>
<GID>744</GID>
<name>IN_2</name></connection>
<intersection>507.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>507.5,-111.5,507.5,-77</points>
<intersection>-111.5 5</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-111.5,507.5,-111.5</points>
<connection>
<GID>689</GID>
<name>OUT_7</name></connection>
<intersection>507.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>508,-88,534,-88</points>
<connection>
<GID>728</GID>
<name>IN_2</name></connection>
<connection>
<GID>745</GID>
<name>IN_2</name></connection>
<intersection>508 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>508,-112.5,508,-88</points>
<intersection>-112.5 5</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-112.5,508,-112.5</points>
<connection>
<GID>689</GID>
<name>OUT_6</name></connection>
<intersection>508 4</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-109.5,497,-73</points>
<intersection>-109.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-73,497,-73</points>
<connection>
<GID>757</GID>
<name>OUT_2</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-109.5,498,-109.5</points>
<connection>
<GID>689</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>508.5,-99,534,-99</points>
<connection>
<GID>729</GID>
<name>IN_2</name></connection>
<connection>
<GID>746</GID>
<name>IN_2</name></connection>
<intersection>508.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>508.5,-113.5,508.5,-99</points>
<intersection>-113.5 7</intersection>
<intersection>-99 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>503,-113.5,508.5,-113.5</points>
<connection>
<GID>689</GID>
<name>OUT_5</name></connection>
<intersection>508.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-122.5,497,-72</points>
<intersection>-122.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>487,-72,497,-72</points>
<connection>
<GID>757</GID>
<name>OUT_3</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,-122.5,498,-122.5</points>
<connection>
<GID>687</GID>
<name>load</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509,-108.5,534,-108.5</points>
<connection>
<GID>730</GID>
<name>IN_2</name></connection>
<connection>
<GID>747</GID>
<name>IN_2</name></connection>
<intersection>509 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>509,-114.5,509,-108.5</points>
<intersection>-114.5 5</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-114.5,509,-114.5</points>
<connection>
<GID>689</GID>
<name>OUT_4</name></connection>
<intersection>509 4</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485.5,-95,485.5,-78</points>
<intersection>-95 2</intersection>
<intersection>-87 8</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480.5,-78,485.5,-78</points>
<intersection>480.5 3</intersection>
<intersection>485.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>472,-95,485.5,-95</points>
<intersection>472 5</intersection>
<intersection>485.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>480.5,-78,480.5,-74</points>
<intersection>-78 1</intersection>
<intersection>-74 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>480.5,-74,481,-74</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<intersection>480.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>472,-109,472,-95</points>
<intersection>-109 6</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>439,-109,472,-109</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<intersection>472 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>483.5,-87,485.5,-87</points>
<connection>
<GID>760</GID>
<name>OUT_1</name></connection>
<intersection>485.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509.5,-119.5,534,-119.5</points>
<connection>
<GID>731</GID>
<name>IN_2</name></connection>
<connection>
<GID>748</GID>
<name>IN_2</name></connection>
<intersection>509.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>509.5,-119.5,509.5,-115.5</points>
<intersection>-119.5 1</intersection>
<intersection>-115.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-115.5,509.5,-115.5</points>
<connection>
<GID>689</GID>
<name>OUT_3</name></connection>
<intersection>509.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>486,-95.5,486,-78.5</points>
<intersection>-95.5 2</intersection>
<intersection>-89 8</intersection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>480,-78.5,486,-78.5</points>
<intersection>480 3</intersection>
<intersection>486 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>472.5,-95.5,486,-95.5</points>
<intersection>472.5 5</intersection>
<intersection>486 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>480,-78.5,480,-75</points>
<intersection>-78.5 1</intersection>
<intersection>-75 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>480,-75,481,-75</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>480 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>472.5,-110,472.5,-95.5</points>
<intersection>-110 6</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>439,-110,472.5,-110</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>472.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>483.5,-89,486,-89</points>
<connection>
<GID>760</GID>
<name>OUT_0</name></connection>
<intersection>486 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>510,-130.5,534,-130.5</points>
<connection>
<GID>732</GID>
<name>IN_2</name></connection>
<connection>
<GID>749</GID>
<name>IN_2</name></connection>
<intersection>510 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>510,-130.5,510,-116.5</points>
<intersection>-130.5 1</intersection>
<intersection>-116.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-116.5,510,-116.5</points>
<connection>
<GID>689</GID>
<name>OUT_2</name></connection>
<intersection>510 4</intersection></hsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>510.5,-141,534,-141</points>
<connection>
<GID>733</GID>
<name>IN_2</name></connection>
<connection>
<GID>750</GID>
<name>IN_2</name></connection>
<intersection>510.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>510.5,-141,510.5,-117.5</points>
<intersection>-141 2</intersection>
<intersection>-117.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-117.5,510.5,-117.5</points>
<connection>
<GID>689</GID>
<name>OUT_1</name></connection>
<intersection>510.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>511,-152,534,-152</points>
<connection>
<GID>734</GID>
<name>IN_2</name></connection>
<connection>
<GID>751</GID>
<name>IN_2</name></connection>
<intersection>511 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>511,-152,511,-118.5</points>
<intersection>-152 1</intersection>
<intersection>-118.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-118.5,511,-118.5</points>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection>
<intersection>511 4</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>511.5,-79,534,-79</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<connection>
<GID>744</GID>
<name>IN_1</name></connection>
<intersection>511.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>511.5,-98,511.5,-79</points>
<intersection>-98 5</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-98,511.5,-98</points>
<connection>
<GID>725</GID>
<name>OUT_7</name></connection>
<intersection>511.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>512,-90,534,-90</points>
<connection>
<GID>728</GID>
<name>IN_1</name></connection>
<connection>
<GID>745</GID>
<name>IN_1</name></connection>
<intersection>512 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>512,-99,512,-90</points>
<intersection>-99 5</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-99,512,-99</points>
<connection>
<GID>725</GID>
<name>OUT_6</name></connection>
<intersection>512 4</intersection></hsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503,-100,534,-100</points>
<connection>
<GID>725</GID>
<name>OUT_5</name></connection>
<intersection>521.5 9</intersection>
<intersection>534 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>534,-101,534,-100</points>
<connection>
<GID>746</GID>
<name>IN_1</name></connection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>521.5,-101,521.5,-100</points>
<connection>
<GID>729</GID>
<name>IN_1</name></connection>
<intersection>-100 1</intersection></vsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>513,-110.5,534,-110.5</points>
<connection>
<GID>730</GID>
<name>IN_1</name></connection>
<connection>
<GID>747</GID>
<name>IN_1</name></connection>
<intersection>513 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>513,-110.5,513,-101</points>
<intersection>-110.5 1</intersection>
<intersection>-101 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-101,513,-101</points>
<connection>
<GID>725</GID>
<name>OUT_4</name></connection>
<intersection>513 4</intersection></hsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>513.5,-121.5,534,-121.5</points>
<connection>
<GID>731</GID>
<name>IN_1</name></connection>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>513.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>513.5,-121.5,513.5,-102</points>
<intersection>-121.5 1</intersection>
<intersection>-102 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-102,513.5,-102</points>
<connection>
<GID>725</GID>
<name>OUT_3</name></connection>
<intersection>513.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>514,-132.5,534,-132.5</points>
<connection>
<GID>732</GID>
<name>IN_1</name></connection>
<connection>
<GID>749</GID>
<name>IN_1</name></connection>
<intersection>514 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>514,-132.5,514,-103</points>
<intersection>-132.5 1</intersection>
<intersection>-103 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503,-103,514,-103</points>
<connection>
<GID>725</GID>
<name>OUT_2</name></connection>
<intersection>514 4</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>384.503,1530.65,1020.62,1194.7</PageViewport>
<gate>
<ID>1497</ID>
<type>AA_LABEL</type>
<position>652.5,1381.5</position>
<gparam>LABEL_TEXT Skip to page 9</gparam>
<gparam>TEXT_HEIGHT 20</gparam>
<gparam>angle 0.0</gparam></gate></page 7>
<page 8>
<PageViewport>386.325,1442.33,759.325,1245.34</PageViewport>
<gate>
<ID>1538</ID>
<type>DA_FROM</type>
<position>405,1338.5</position>
<input>
<ID>IN_0</ID>2073 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>1540</ID>
<type>DE_TO</type>
<position>415,1340.5</position>
<input>
<ID>IN_0</ID>2074 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WE</lparam></gate>
<gate>
<ID>1541</ID>
<type>DA_FROM</type>
<position>426.5,1371.5</position>
<input>
<ID>IN_0</ID>2076 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LD/ST</lparam></gate>
<gate>
<ID>1543</ID>
<type>AA_LABEL</type>
<position>446.5,1386.5</position>
<gparam>LABEL_TEXT MAR-in</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1545</ID>
<type>AA_LABEL</type>
<position>497.5,1418</position>
<gparam>LABEL_TEXT Manually</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1547</ID>
<type>AE_SMALL_INVERTER</type>
<position>548,1394.5</position>
<input>
<ID>IN_0</ID>1632 </input>
<output>
<ID>OUT_0</ID>2080 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1549</ID>
<type>BE_NOR2</type>
<position>725.5,1302.5</position>
<input>
<ID>IN_0</ID>2041 </input>
<input>
<ID>IN_1</ID>1465 </input>
<output>
<ID>OUT</ID>2091 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1551</ID>
<type>DE_TO</type>
<position>667.5,1352.5</position>
<input>
<ID>IN_0</ID>2092 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD(0/1)</lparam></gate>
<gate>
<ID>1553</ID>
<type>DE_TO</type>
<position>667.5,1365.5</position>
<input>
<ID>IN_0</ID>2093 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ST(0/1)</lparam></gate>
<gate>
<ID>1555</ID>
<type>DA_FROM</type>
<position>400,1327.5</position>
<input>
<ID>IN_0</ID>2094 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ST(0/1)</lparam></gate>
<gate>
<ID>1557</ID>
<type>DA_FROM</type>
<position>423,1308</position>
<input>
<ID>IN_0</ID>2095 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD(0/1)</lparam></gate>
<gate>
<ID>1559</ID>
<type>DE_TO</type>
<position>451,1279</position>
<input>
<ID>IN_0</ID>1762 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1561</ID>
<type>DA_FROM</type>
<position>538.5,1373</position>
<input>
<ID>IN_0</ID>2096 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1563</ID>
<type>DA_FROM</type>
<position>569.5,1379.5</position>
<input>
<ID>IN_0</ID>2097 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1565</ID>
<type>DA_FROM</type>
<position>592,1388.5</position>
<input>
<ID>IN_0</ID>2098 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1567</ID>
<type>DA_FROM</type>
<position>607,1340</position>
<input>
<ID>IN_0</ID>2099 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1569</ID>
<type>DA_FROM</type>
<position>723,1288.5</position>
<input>
<ID>IN_0</ID>2100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>1573</ID>
<type>EE_VDD</type>
<position>534,1394</position>
<output>
<ID>OUT_0</ID>2102 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>841</ID>
<type>EE_VDD</type>
<position>710.5,1298.5</position>
<output>
<ID>OUT_0</ID>1028 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>846</ID>
<type>DA_FROM</type>
<position>678.5,1305.5</position>
<input>
<ID>IN_0</ID>1464 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr0</lparam></gate>
<gate>
<ID>847</ID>
<type>AE_OR2</type>
<position>668,1361</position>
<input>
<ID>IN_0</ID>2093 </input>
<input>
<ID>IN_1</ID>1625 </input>
<output>
<ID>OUT</ID>1027 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>964</ID>
<type>DA_FROM</type>
<position>678.5,1307.5</position>
<input>
<ID>IN_0</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr1</lparam></gate>
<gate>
<ID>965</ID>
<type>AE_OR2</type>
<position>668,1357</position>
<input>
<ID>IN_0</ID>2092 </input>
<input>
<ID>IN_1</ID>1554 </input>
<output>
<ID>OUT</ID>834 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>966</ID>
<type>DA_FROM</type>
<position>678.5,1309.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr2</lparam></gate>
<gate>
<ID>967</ID>
<type>DE_TO</type>
<position>673.5,1357</position>
<input>
<ID>IN_0</ID>834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD</lparam></gate>
<gate>
<ID>968</ID>
<type>DA_FROM</type>
<position>678.5,1311.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr3</lparam></gate>
<gate>
<ID>969</ID>
<type>DE_TO</type>
<position>673.5,1361</position>
<input>
<ID>IN_0</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>970</ID>
<type>DA_FROM</type>
<position>678.5,1313.5</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr4</lparam></gate>
<gate>
<ID>971</ID>
<type>DA_FROM</type>
<position>678.5,1315.5</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr5</lparam></gate>
<gate>
<ID>972</ID>
<type>DA_FROM</type>
<position>678.5,1317.5</position>
<input>
<ID>IN_0</ID>1206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr6</lparam></gate>
<gate>
<ID>973</ID>
<type>DE_TO</type>
<position>661,1344</position>
<input>
<ID>IN_0</ID>1029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>975</ID>
<type>DA_FROM</type>
<position>678.5,1319.5</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr7</lparam></gate>
<gate>
<ID>976</ID>
<type>DE_TO</type>
<position>661,1338.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>977</ID>
<type>AA_LABEL</type>
<position>513,1400.5</position>
<gparam>LABEL_TEXT Enter with keypads</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>988</ID>
<type>AA_LABEL</type>
<position>628,1410</position>
<gparam>LABEL_TEXT Offset decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>990</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>694,1308</position>
<input>
<ID>ENABLE_0</ID>1465 </input>
<input>
<ID>IN_1</ID>1464 </input>
<input>
<ID>IN_11</ID>1035 </input>
<input>
<ID>IN_13</ID>1206 </input>
<input>
<ID>IN_15</ID>1056 </input>
<input>
<ID>IN_3</ID>1042 </input>
<input>
<ID>IN_5</ID>1173 </input>
<input>
<ID>IN_7</ID>1031 </input>
<input>
<ID>IN_9</ID>1034 </input>
<output>
<ID>OUT_1</ID>2040 </output>
<output>
<ID>OUT_11</ID>2034 </output>
<output>
<ID>OUT_13</ID>2036 </output>
<output>
<ID>OUT_15</ID>2033 </output>
<output>
<ID>OUT_3</ID>2039 </output>
<output>
<ID>OUT_5</ID>2038 </output>
<output>
<ID>OUT_7</ID>2035 </output>
<output>
<ID>OUT_9</ID>2037 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>993</ID>
<type>DA_FROM</type>
<position>689.5,1317.5</position>
<input>
<ID>IN_0</ID>1465 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD</lparam></gate>
<gate>
<ID>994</ID>
<type>AA_LABEL</type>
<position>714,1301.5</position>
<gparam>LABEL_TEXT CC decoder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>996</ID>
<type>AA_LABEL</type>
<position>741,1295</position>
<gparam>LABEL_TEXT CC Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1000</ID>
<type>AA_LABEL</type>
<position>746,1326</position>
<gparam>LABEL_TEXT Do we branch?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1002</ID>
<type>DA_FROM</type>
<position>430,1344</position>
<input>
<ID>IN_0</ID>1044 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WE</lparam></gate>
<gate>
<ID>1005</ID>
<type>DA_FROM</type>
<position>527,1338</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr0</lparam></gate>
<gate>
<ID>1006</ID>
<type>DA_FROM</type>
<position>527,1340</position>
<input>
<ID>IN_0</ID>1150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr1</lparam></gate>
<gate>
<ID>1007</ID>
<type>DA_FROM</type>
<position>527,1342</position>
<input>
<ID>IN_0</ID>1145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr2</lparam></gate>
<gate>
<ID>1008</ID>
<type>DA_FROM</type>
<position>527,1344</position>
<input>
<ID>IN_0</ID>1083 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr3</lparam></gate>
<gate>
<ID>1009</ID>
<type>DA_FROM</type>
<position>527,1346</position>
<input>
<ID>IN_0</ID>1082 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr4</lparam></gate>
<gate>
<ID>1011</ID>
<type>DA_FROM</type>
<position>527,1348</position>
<input>
<ID>IN_0</ID>1079 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr5</lparam></gate>
<gate>
<ID>1013</ID>
<type>DA_FROM</type>
<position>527,1350</position>
<input>
<ID>IN_0</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr6</lparam></gate>
<gate>
<ID>1014</ID>
<type>DA_FROM</type>
<position>527,1352</position>
<input>
<ID>IN_0</ID>1061 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr7</lparam></gate>
<gate>
<ID>1015</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>560,1348.5</position>
<input>
<ID>ENABLE_0</ID>1995 </input>
<input>
<ID>IN_0</ID>1057 </input>
<input>
<ID>IN_1</ID>1150 </input>
<input>
<ID>IN_2</ID>1145 </input>
<input>
<ID>IN_3</ID>1083 </input>
<input>
<ID>IN_4</ID>1082 </input>
<input>
<ID>IN_5</ID>1079 </input>
<input>
<ID>IN_6</ID>1078 </input>
<input>
<ID>IN_7</ID>1061 </input>
<output>
<ID>OUT_0</ID>1974 </output>
<output>
<ID>OUT_1</ID>1971 </output>
<output>
<ID>OUT_2</ID>1992 </output>
<output>
<ID>OUT_3</ID>1970 </output>
<output>
<ID>OUT_4</ID>1973 </output>
<output>
<ID>OUT_5</ID>1993 </output>
<output>
<ID>OUT_6</ID>1972 </output>
<output>
<ID>OUT_7</ID>1994 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1022</ID>
<type>AA_AND2</type>
<position>737,1321.5</position>
<input>
<ID>IN_0</ID>1964 </input>
<input>
<ID>IN_1</ID>1611 </input>
<output>
<ID>OUT</ID>1499 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1026</ID>
<type>AA_AND2</type>
<position>737,1317.5</position>
<input>
<ID>IN_0</ID>1969 </input>
<input>
<ID>IN_1</ID>1610 </input>
<output>
<ID>OUT</ID>1493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1028</ID>
<type>AA_AND2</type>
<position>737,1313.5</position>
<input>
<ID>IN_0</ID>1612 </input>
<input>
<ID>IN_1</ID>1607 </input>
<output>
<ID>OUT</ID>1470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1033</ID>
<type>AE_OR3</type>
<position>743.5,1317.5</position>
<input>
<ID>IN_0</ID>1499 </input>
<input>
<ID>IN_1</ID>1493 </input>
<input>
<ID>IN_2</ID>1470 </input>
<output>
<ID>OUT</ID>1500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1035</ID>
<type>AA_AND2</type>
<position>751,1318.5</position>
<input>
<ID>IN_0</ID>1501 </input>
<input>
<ID>IN_1</ID>1500 </input>
<output>
<ID>OUT</ID>1515 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1052</ID>
<type>AA_AND2</type>
<position>656,1338.5</position>
<input>
<ID>IN_0</ID>1594 </input>
<input>
<ID>IN_1</ID>1555 </input>
<output>
<ID>OUT</ID>1030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1053</ID>
<type>AA_AND2</type>
<position>656,1333</position>
<input>
<ID>IN_0</ID>1594 </input>
<input>
<ID>IN_1</ID>1606 </input>
<output>
<ID>OUT</ID>1947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1054</ID>
<type>BE_NOR2</type>
<position>644.5,1353</position>
<input>
<ID>IN_0</ID>1594 </input>
<input>
<ID>IN_1</ID>1606 </input>
<output>
<ID>OUT</ID>1951 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1055</ID>
<type>BA_DECODER_2x4</type>
<position>660.5,1359</position>
<input>
<ID>ENABLE</ID>1951 </input>
<input>
<ID>IN_0</ID>1969 </input>
<input>
<ID>IN_1</ID>1964 </input>
<output>
<ID>OUT_0</ID>1554 </output>
<output>
<ID>OUT_1</ID>2092 </output>
<output>
<ID>OUT_2</ID>1625 </output>
<output>
<ID>OUT_3</ID>2093 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1056</ID>
<type>DA_FROM</type>
<position>746,1322.5</position>
<input>
<ID>IN_0</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRop</lparam></gate>
<gate>
<ID>1057</ID>
<type>AA_LABEL</type>
<position>655.5,1341.5</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1058</ID>
<type>AA_LABEL</type>
<position>655.5,1347</position>
<gparam>LABEL_TEXT ADD</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1059</ID>
<type>AA_LABEL</type>
<position>656,1336</position>
<gparam>LABEL_TEXT BRnzp</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1060</ID>
<type>DM_NOR8</type>
<position>707,1290.5</position>
<input>
<ID>IN_0</ID>2033 </input>
<input>
<ID>IN_1</ID>2036 </input>
<input>
<ID>IN_2</ID>2034 </input>
<input>
<ID>IN_3</ID>2037 </input>
<input>
<ID>IN_4</ID>2040 </input>
<input>
<ID>IN_5</ID>2039 </input>
<input>
<ID>IN_6</ID>2038 </input>
<input>
<ID>IN_7</ID>2035 </input>
<output>
<ID>OUT</ID>1595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1061</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>521,1395</position>
<input>
<ID>ENABLE_0</ID>1568 </input>
<input>
<ID>IN_0</ID>1569 </input>
<input>
<ID>IN_1</ID>1570 </input>
<input>
<ID>IN_2</ID>1571 </input>
<input>
<ID>IN_3</ID>1572 </input>
<input>
<ID>IN_4</ID>1573 </input>
<input>
<ID>IN_5</ID>1574 </input>
<input>
<ID>IN_6</ID>1575 </input>
<input>
<ID>IN_7</ID>1576 </input>
<output>
<ID>OUT_0</ID>1557 </output>
<output>
<ID>OUT_1</ID>1558 </output>
<output>
<ID>OUT_2</ID>1559 </output>
<output>
<ID>OUT_3</ID>1560 </output>
<output>
<ID>OUT_4</ID>1561 </output>
<output>
<ID>OUT_5</ID>1562 </output>
<output>
<ID>OUT_6</ID>1563 </output>
<output>
<ID>OUT_7</ID>1564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1063</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>521,1383</position>
<input>
<ID>ENABLE_0</ID>1567 </input>
<input>
<ID>IN_0</ID>2055 </input>
<input>
<ID>IN_1</ID>2057 </input>
<input>
<ID>IN_2</ID>2053 </input>
<input>
<ID>IN_3</ID>2058 </input>
<input>
<ID>IN_4</ID>2054 </input>
<input>
<ID>IN_5</ID>2056 </input>
<input>
<ID>IN_6</ID>2059 </input>
<input>
<ID>IN_7</ID>2060 </input>
<output>
<ID>OUT_0</ID>1557 </output>
<output>
<ID>OUT_1</ID>1558 </output>
<output>
<ID>OUT_2</ID>1559 </output>
<output>
<ID>OUT_3</ID>1560 </output>
<output>
<ID>OUT_4</ID>1561 </output>
<output>
<ID>OUT_5</ID>1562 </output>
<output>
<ID>OUT_6</ID>1563 </output>
<output>
<ID>OUT_7</ID>1564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1065</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>534,1387</position>
<input>
<ID>ENABLE_0</ID>2102 </input>
<input>
<ID>IN_0</ID>1557 </input>
<input>
<ID>IN_1</ID>1558 </input>
<input>
<ID>IN_2</ID>1559 </input>
<input>
<ID>IN_3</ID>1560 </input>
<input>
<ID>IN_4</ID>1561 </input>
<input>
<ID>IN_5</ID>1562 </input>
<input>
<ID>IN_6</ID>1563 </input>
<input>
<ID>IN_7</ID>1564 </input>
<output>
<ID>OUT_0</ID>1579 </output>
<output>
<ID>OUT_1</ID>1582 </output>
<output>
<ID>OUT_2</ID>1583 </output>
<output>
<ID>OUT_3</ID>1581 </output>
<output>
<ID>OUT_4</ID>1584 </output>
<output>
<ID>OUT_5</ID>1578 </output>
<output>
<ID>OUT_6</ID>1577 </output>
<output>
<ID>OUT_7</ID>1580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1067</ID>
<type>BA_DECODER_2x4</type>
<position>516,1404</position>
<input>
<ID>ENABLE</ID>1565 </input>
<input>
<ID>IN_0</ID>1566 </input>
<output>
<ID>OUT_0</ID>1567 </output>
<output>
<ID>OUT_1</ID>1568 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1069</ID>
<type>EE_VDD</type>
<position>513,1408</position>
<output>
<ID>OUT_0</ID>1565 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1071</ID>
<type>AE_SMALL_INVERTER</type>
<position>651,1341</position>
<input>
<ID>IN_0</ID>1606 </input>
<output>
<ID>OUT_0</ID>1555 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1072</ID>
<type>AA_TOGGLE</type>
<position>510.5,1402.5</position>
<output>
<ID>OUT_0</ID>1566 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1073</ID>
<type>DD_KEYPAD_HEX</type>
<position>498,1409.5</position>
<output>
<ID>OUT_0</ID>1573 </output>
<output>
<ID>OUT_1</ID>1574 </output>
<output>
<ID>OUT_2</ID>1575 </output>
<output>
<ID>OUT_3</ID>1576 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>1074</ID>
<type>DD_KEYPAD_HEX</type>
<position>498,1397</position>
<output>
<ID>OUT_0</ID>1569 </output>
<output>
<ID>OUT_1</ID>1570 </output>
<output>
<ID>OUT_2</ID>1571 </output>
<output>
<ID>OUT_3</ID>1572 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>1075</ID>
<type>BA_DECODER_2x4</type>
<position>714.5,1294.5</position>
<input>
<ID>ENABLE</ID>1028 </input>
<input>
<ID>IN_0</ID>1595 </input>
<input>
<ID>IN_1</ID>2033 </input>
<output>
<ID>OUT_0</ID>1607 </output>
<output>
<ID>OUT_1</ID>1610 </output>
<output>
<ID>OUT_2</ID>1611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1077</ID>
<type>AE_SMALL_INVERTER</type>
<position>651,1345</position>
<input>
<ID>IN_0</ID>1594 </input>
<output>
<ID>OUT_0</ID>1605 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1080</ID>
<type>AA_LABEL</type>
<position>719,1294</position>
<gparam>LABEL_TEXT nzp</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>1081</ID>
<type>AA_LABEL</type>
<position>608,1383</position>
<gparam>LABEL_TEXT Always Write or Output</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1082</ID>
<type>EE_VDD</type>
<position>572.5,1300.5</position>
<output>
<ID>OUT_0</ID>1617 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1083</ID>
<type>EE_VDD</type>
<position>572.5,1323.5</position>
<output>
<ID>OUT_0</ID>1618 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1084</ID>
<type>AA_REGISTER4</type>
<position>726.5,1294</position>
<input>
<ID>IN_0</ID>1607 </input>
<input>
<ID>IN_1</ID>1610 </input>
<input>
<ID>IN_2</ID>1611 </input>
<input>
<ID>clock</ID>2100 </input>
<input>
<ID>load</ID>2091 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1089</ID>
<type>AA_LABEL</type>
<position>415.5,1322.5</position>
<gparam>LABEL_TEXT Bits 0-1</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1090</ID>
<type>AA_LABEL</type>
<position>415.5,1325</position>
<gparam>LABEL_TEXT Bits 2-3</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1091</ID>
<type>AA_LABEL</type>
<position>416,1321.5</position>
<gparam>LABEL_TEXT Read output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1092</ID>
<type>AA_LABEL</type>
<position>416,1326.5</position>
<gparam>LABEL_TEXT Read output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1094</ID>
<type>AA_LABEL</type>
<position>579,1343.5</position>
<gparam>LABEL_TEXT Input tri-bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1095</ID>
<type>AA_AND2</type>
<position>605.5,1322.5</position>
<input>
<ID>IN_0</ID>1696 </input>
<input>
<ID>IN_1</ID>1695 </input>
<output>
<ID>OUT</ID>1714 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1096</ID>
<type>AA_LABEL</type>
<position>423.5,1304.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1097</ID>
<type>AA_LABEL</type>
<position>424,1303</position>
<gparam>LABEL_TEXT R0-R3</gparam>
<gparam>TEXT_HEIGHT 0.75</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1098</ID>
<type>AA_AND2</type>
<position>600.5,1326</position>
<input>
<ID>IN_0</ID>1698 </input>
<input>
<ID>IN_1</ID>1697 </input>
<output>
<ID>OUT</ID>1715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1099</ID>
<type>AA_LABEL</type>
<position>517.5,1373</position>
<gparam>LABEL_TEXT ClockOn-LoadOff  = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1100</ID>
<type>AA_LABEL</type>
<position>517.5,1371.5</position>
<gparam>LABEL_TEXT ClockOff-LoadOn  = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1101</ID>
<type>AA_AND2</type>
<position>605.5,1329.5</position>
<input>
<ID>IN_0</ID>1700 </input>
<input>
<ID>IN_1</ID>1699 </input>
<output>
<ID>OUT</ID>1716 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1102</ID>
<type>AE_REGISTER8</type>
<position>549,1386.5</position>
<input>
<ID>IN_0</ID>1579 </input>
<input>
<ID>IN_1</ID>1582 </input>
<input>
<ID>IN_2</ID>1583 </input>
<input>
<ID>IN_3</ID>1581 </input>
<input>
<ID>IN_4</ID>1584 </input>
<input>
<ID>IN_5</ID>1578 </input>
<input>
<ID>IN_6</ID>1577 </input>
<input>
<ID>IN_7</ID>1580 </input>
<output>
<ID>OUT_0</ID>1838 </output>
<output>
<ID>OUT_1</ID>1968 </output>
<output>
<ID>OUT_2</ID>1836 </output>
<output>
<ID>OUT_3</ID>1835 </output>
<output>
<ID>OUT_4</ID>1834 </output>
<output>
<ID>OUT_5</ID>1833 </output>
<output>
<ID>OUT_6</ID>1832 </output>
<output>
<ID>OUT_7</ID>1831 </output>
<input>
<ID>clear</ID>1644 </input>
<input>
<ID>clock</ID>2075 </input>
<input>
<ID>count_enable</ID>1632 </input>
<input>
<ID>count_up</ID>1632 </input>
<input>
<ID>load</ID>2080 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 134</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1103</ID>
<type>AE_REGISTER8</type>
<position>450,1287.5</position>
<input>
<ID>IN_0</ID>1782 </input>
<input>
<ID>IN_1</ID>1781 </input>
<input>
<ID>IN_2</ID>1780 </input>
<input>
<ID>IN_3</ID>1779 </input>
<input>
<ID>IN_4</ID>1778 </input>
<input>
<ID>IN_5</ID>1777 </input>
<input>
<ID>IN_6</ID>1776 </input>
<input>
<ID>IN_7</ID>1775 </input>
<output>
<ID>OUT_0</ID>1730 </output>
<output>
<ID>OUT_1</ID>1729 </output>
<output>
<ID>OUT_2</ID>1556 </output>
<output>
<ID>OUT_3</ID>1728 </output>
<output>
<ID>OUT_4</ID>1727 </output>
<output>
<ID>OUT_5</ID>1726 </output>
<output>
<ID>OUT_6</ID>1725 </output>
<output>
<ID>OUT_7</ID>1785 </output>
<input>
<ID>clock</ID>1762 </input>
<input>
<ID>load</ID>1599 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 88</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1104</ID>
<type>AE_REGISTER8</type>
<position>570.5,1386.5</position>
<input>
<ID>IN_0</ID>1868 </input>
<input>
<ID>IN_1</ID>1869 </input>
<input>
<ID>IN_2</ID>1870 </input>
<input>
<ID>IN_3</ID>1871 </input>
<input>
<ID>IN_4</ID>1872 </input>
<input>
<ID>IN_5</ID>1873 </input>
<input>
<ID>IN_6</ID>1867 </input>
<input>
<ID>IN_7</ID>1866 </input>
<output>
<ID>OUT_0</ID>1634 </output>
<output>
<ID>OUT_1</ID>1633 </output>
<output>
<ID>OUT_2</ID>1631 </output>
<output>
<ID>OUT_3</ID>1630 </output>
<output>
<ID>OUT_4</ID>1629 </output>
<output>
<ID>OUT_5</ID>1628 </output>
<output>
<ID>OUT_6</ID>1627 </output>
<output>
<ID>OUT_7</ID>1626 </output>
<input>
<ID>clear</ID>1644 </input>
<input>
<ID>clock</ID>2097 </input>
<input>
<ID>load</ID>1874 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 138</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1105</ID>
<type>AE_REGISTER8</type>
<position>450,1300.5</position>
<input>
<ID>IN_0</ID>1782 </input>
<input>
<ID>IN_1</ID>1781 </input>
<input>
<ID>IN_2</ID>1780 </input>
<input>
<ID>IN_3</ID>1779 </input>
<input>
<ID>IN_4</ID>1778 </input>
<input>
<ID>IN_5</ID>1777 </input>
<input>
<ID>IN_6</ID>1776 </input>
<input>
<ID>IN_7</ID>1775 </input>
<output>
<ID>OUT_0</ID>1738 </output>
<output>
<ID>OUT_1</ID>1737 </output>
<output>
<ID>OUT_2</ID>1736 </output>
<output>
<ID>OUT_3</ID>1735 </output>
<output>
<ID>OUT_4</ID>1734 </output>
<output>
<ID>OUT_5</ID>1733 </output>
<output>
<ID>OUT_6</ID>1732 </output>
<output>
<ID>OUT_7</ID>1731 </output>
<input>
<ID>clock</ID>1762 </input>
<input>
<ID>load</ID>1598 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1106</ID>
<type>AE_REGISTER8</type>
<position>608,1348</position>
<input>
<ID>IN_0</ID>1654 </input>
<input>
<ID>IN_1</ID>1655 </input>
<input>
<ID>IN_2</ID>1656 </input>
<input>
<ID>IN_3</ID>1657 </input>
<input>
<ID>IN_4</ID>1658 </input>
<input>
<ID>IN_5</ID>1653 </input>
<input>
<ID>IN_6</ID>1660 </input>
<input>
<ID>IN_7</ID>1659 </input>
<output>
<ID>OUT_0</ID>1642 </output>
<output>
<ID>OUT_1</ID>1641 </output>
<output>
<ID>OUT_2</ID>1640 </output>
<output>
<ID>OUT_3</ID>1639 </output>
<output>
<ID>OUT_4</ID>1638 </output>
<output>
<ID>OUT_5</ID>1637 </output>
<output>
<ID>OUT_6</ID>1636 </output>
<output>
<ID>OUT_7</ID>1635 </output>
<input>
<ID>clear</ID>1644 </input>
<input>
<ID>clock</ID>2099 </input>
<input>
<ID>load</ID>2072 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1107</ID>
<type>AE_RAM_8x8</type>
<position>585,1387</position>
<input>
<ID>ADDRESS_0</ID>1634 </input>
<input>
<ID>ADDRESS_1</ID>1633 </input>
<input>
<ID>ADDRESS_2</ID>1631 </input>
<input>
<ID>ADDRESS_3</ID>1630 </input>
<input>
<ID>ADDRESS_4</ID>1629 </input>
<input>
<ID>ADDRESS_5</ID>1628 </input>
<input>
<ID>ADDRESS_6</ID>1627 </input>
<input>
<ID>ADDRESS_7</ID>1626 </input>
<input>
<ID>DATA_IN_0</ID>1661 </input>
<input>
<ID>DATA_IN_1</ID>1646 </input>
<input>
<ID>DATA_IN_2</ID>1647 </input>
<input>
<ID>DATA_IN_3</ID>1648 </input>
<input>
<ID>DATA_IN_4</ID>1649 </input>
<input>
<ID>DATA_IN_5</ID>1650 </input>
<input>
<ID>DATA_IN_6</ID>1651 </input>
<input>
<ID>DATA_IN_7</ID>1652 </input>
<output>
<ID>DATA_OUT_0</ID>1661 </output>
<output>
<ID>DATA_OUT_1</ID>1646 </output>
<output>
<ID>DATA_OUT_2</ID>1647 </output>
<output>
<ID>DATA_OUT_3</ID>1648 </output>
<output>
<ID>DATA_OUT_4</ID>1649 </output>
<output>
<ID>DATA_OUT_5</ID>1650 </output>
<output>
<ID>DATA_OUT_6</ID>1651 </output>
<output>
<ID>DATA_OUT_7</ID>1652 </output>
<input>
<ID>ENABLE_0</ID>1786 </input>
<input>
<ID>write_clock</ID>2098 </input>
<input>
<ID>write_enable</ID>1645 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:13 83</lparam>
<lparam>Address:14 83</lparam>
<lparam>Address:15 83</lparam>
<lparam>Address:16 83</lparam>
<lparam>Address:17 83</lparam>
<lparam>Address:23 46</lparam>
<lparam>Address:24 71</lparam>
<lparam>Address:25 135</lparam>
<lparam>Address:26 1</lparam>
<lparam>Address:28 36</lparam>
<lparam>Address:56 1</lparam>
<lparam>Address:58 255</lparam>
<lparam>Address:81 4</lparam>
<lparam>Address:83 13</lparam>
<lparam>Address:84 2</lparam>
<lparam>Address:87 221</lparam>
<lparam>Address:88 46</lparam>
<lparam>Address:133 250</lparam>
<lparam>Address:138 52</lparam></gate>
<gate>
<ID>1108</ID>
<type>AE_REGISTER8</type>
<position>625.5,1348</position>
<input>
<ID>IN_0</ID>2064 </input>
<input>
<ID>IN_1</ID>2068 </input>
<input>
<ID>IN_2</ID>2067 </input>
<input>
<ID>IN_3</ID>2065 </input>
<input>
<ID>IN_4</ID>2063 </input>
<input>
<ID>IN_5</ID>2066 </input>
<input>
<ID>IN_6</ID>2069 </input>
<input>
<ID>IN_7</ID>2062 </input>
<output>
<ID>OUT_0</ID>1616 </output>
<output>
<ID>OUT_1</ID>1614 </output>
<output>
<ID>OUT_2</ID>1613 </output>
<output>
<ID>OUT_3</ID>1612 </output>
<output>
<ID>OUT_4</ID>1969 </output>
<output>
<ID>OUT_5</ID>1964 </output>
<output>
<ID>OUT_6</ID>1606 </output>
<output>
<ID>OUT_7</ID>1594 </output>
<input>
<ID>clear</ID>1644 </input>
<input>
<ID>clock</ID>2099 </input>
<input>
<ID>load</ID>2088 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1109</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>411,1277.5</position>
<input>
<ID>ENABLE_0</ID>2002 </input>
<input>
<ID>IN_0</ID>1984 </input>
<input>
<ID>IN_1</ID>1991 </input>
<input>
<ID>IN_2</ID>1990 </input>
<input>
<ID>IN_3</ID>1989 </input>
<input>
<ID>IN_4</ID>1988 </input>
<input>
<ID>IN_5</ID>1987 </input>
<input>
<ID>IN_6</ID>1986 </input>
<input>
<ID>IN_7</ID>1985 </input>
<output>
<ID>OUT_0</ID>1782 </output>
<output>
<ID>OUT_1</ID>1781 </output>
<output>
<ID>OUT_2</ID>1780 </output>
<output>
<ID>OUT_3</ID>1779 </output>
<output>
<ID>OUT_4</ID>1778 </output>
<output>
<ID>OUT_5</ID>1777 </output>
<output>
<ID>OUT_6</ID>1776 </output>
<output>
<ID>OUT_7</ID>1775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1110</ID>
<type>BB_CLOCK</type>
<position>444,1279</position>
<output>
<ID>CLK</ID>1762 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1111</ID>
<type>AA_TOGGLE</type>
<position>545,1400.5</position>
<output>
<ID>OUT_0</ID>1632 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1112</ID>
<type>AA_LABEL</type>
<position>498,1416.5</position>
<gparam>LABEL_TEXT load initial address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1113</ID>
<type>AA_LABEL</type>
<position>542.5,1403</position>
<gparam>LABEL_TEXT Count = 1, Don't count = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1114</ID>
<type>AA_TOGGLE</type>
<position>552,1358.5</position>
<output>
<ID>OUT_0</ID>1644 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1115</ID>
<type>AA_LABEL</type>
<position>547,1361</position>
<gparam>LABEL_TEXT Reset Registers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1116</ID>
<type>AA_LABEL</type>
<position>545,1395</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1117</ID>
<type>AA_LABEL</type>
<position>573.5,1396</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1118</ID>
<type>AA_LABEL</type>
<position>585,1395.5</position>
<gparam>LABEL_TEXT RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1119</ID>
<type>AA_LABEL</type>
<position>611.5,1356</position>
<gparam>LABEL_TEXT MDR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1123</ID>
<type>AA_LABEL</type>
<position>599.5,1397.5</position>
<gparam>LABEL_TEXT Write Enable = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1124</ID>
<type>AA_LABEL</type>
<position>599,1395.5</position>
<gparam>LABEL_TEXT Output Enable = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1125</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>591.5,1348.5</position>
<input>
<ID>ENABLE_0</ID>1786 </input>
<input>
<ID>IN_0</ID>1661 </input>
<input>
<ID>IN_1</ID>1646 </input>
<input>
<ID>IN_2</ID>1647 </input>
<input>
<ID>IN_3</ID>1648 </input>
<input>
<ID>IN_4</ID>1649 </input>
<input>
<ID>IN_5</ID>1650 </input>
<input>
<ID>IN_6</ID>1651 </input>
<input>
<ID>IN_7</ID>1652 </input>
<output>
<ID>OUT_0</ID>1654 </output>
<output>
<ID>OUT_1</ID>1655 </output>
<output>
<ID>OUT_2</ID>1656 </output>
<output>
<ID>OUT_3</ID>1657 </output>
<output>
<ID>OUT_4</ID>1658 </output>
<output>
<ID>OUT_5</ID>1653 </output>
<output>
<ID>OUT_6</ID>1660 </output>
<output>
<ID>OUT_7</ID>1659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1126</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>576.5,1348.5</position>
<input>
<ID>ENABLE_0</ID>1645 </input>
<input>
<ID>IN_0</ID>1974 </input>
<input>
<ID>IN_1</ID>1971 </input>
<input>
<ID>IN_2</ID>1992 </input>
<input>
<ID>IN_3</ID>1970 </input>
<input>
<ID>IN_4</ID>1973 </input>
<input>
<ID>IN_5</ID>1993 </input>
<input>
<ID>IN_6</ID>1972 </input>
<input>
<ID>IN_7</ID>1994 </input>
<output>
<ID>OUT_0</ID>1661 </output>
<output>
<ID>OUT_1</ID>1646 </output>
<output>
<ID>OUT_2</ID>1647 </output>
<output>
<ID>OUT_3</ID>1648 </output>
<output>
<ID>OUT_4</ID>1649 </output>
<output>
<ID>OUT_5</ID>1650 </output>
<output>
<ID>OUT_6</ID>1651 </output>
<output>
<ID>OUT_7</ID>1652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1127</ID>
<type>AA_LABEL</type>
<position>626.5,1356</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1128</ID>
<type>AA_LABEL</type>
<position>427,1278.5</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 2.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1129</ID>
<type>AA_AND2</type>
<position>543.5,1374</position>
<input>
<ID>IN_0</ID>1604 </input>
<input>
<ID>IN_1</ID>2096 </input>
<output>
<ID>OUT</ID>2075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1132</ID>
<type>AA_TOGGLE</type>
<position>520.5,1375</position>
<output>
<ID>OUT_0</ID>1604 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1133</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>587.5,1313.5</position>
<input>
<ID>ENABLE_0</ID>1667 </input>
<input>
<ID>IN_0</ID>1822 </input>
<input>
<ID>IN_1</ID>1815 </input>
<input>
<ID>IN_10</ID>1827 </input>
<input>
<ID>IN_11</ID>1828 </input>
<input>
<ID>IN_12</ID>1825 </input>
<input>
<ID>IN_13</ID>1823 </input>
<input>
<ID>IN_14</ID>1826 </input>
<input>
<ID>IN_15</ID>1830 </input>
<input>
<ID>IN_2</ID>1819 </input>
<input>
<ID>IN_3</ID>1818 </input>
<input>
<ID>IN_4</ID>1816 </input>
<input>
<ID>IN_5</ID>1817 </input>
<input>
<ID>IN_6</ID>1820 </input>
<input>
<ID>IN_7</ID>1821 </input>
<input>
<ID>IN_8</ID>1829 </input>
<input>
<ID>IN_9</ID>1824 </input>
<output>
<ID>OUT_0</ID>1685 </output>
<output>
<ID>OUT_1</ID>1686 </output>
<output>
<ID>OUT_10</ID>1695 </output>
<output>
<ID>OUT_11</ID>1696 </output>
<output>
<ID>OUT_12</ID>1697 </output>
<output>
<ID>OUT_13</ID>1698 </output>
<output>
<ID>OUT_14</ID>1699 </output>
<output>
<ID>OUT_15</ID>1700 </output>
<output>
<ID>OUT_2</ID>1687 </output>
<output>
<ID>OUT_3</ID>1688 </output>
<output>
<ID>OUT_4</ID>1689 </output>
<output>
<ID>OUT_5</ID>1690 </output>
<output>
<ID>OUT_6</ID>1691 </output>
<output>
<ID>OUT_7</ID>1692 </output>
<output>
<ID>OUT_8</ID>1693 </output>
<output>
<ID>OUT_9</ID>1694 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1134</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>587.5,1290.5</position>
<input>
<ID>ENABLE_0</ID>1666 </input>
<input>
<ID>IN_0</ID>1799 </input>
<input>
<ID>IN_1</ID>1801 </input>
<input>
<ID>IN_10</ID>1808 </input>
<input>
<ID>IN_11</ID>1810 </input>
<input>
<ID>IN_12</ID>1811 </input>
<input>
<ID>IN_13</ID>1813 </input>
<input>
<ID>IN_14</ID>1812 </input>
<input>
<ID>IN_15</ID>1814 </input>
<input>
<ID>IN_2</ID>1800 </input>
<input>
<ID>IN_3</ID>1802 </input>
<input>
<ID>IN_4</ID>1803 </input>
<input>
<ID>IN_5</ID>1804 </input>
<input>
<ID>IN_6</ID>1806 </input>
<input>
<ID>IN_7</ID>1805 </input>
<input>
<ID>IN_8</ID>1809 </input>
<input>
<ID>IN_9</ID>1807 </input>
<output>
<ID>OUT_0</ID>1669 </output>
<output>
<ID>OUT_1</ID>1677 </output>
<output>
<ID>OUT_10</ID>1674 </output>
<output>
<ID>OUT_11</ID>1682 </output>
<output>
<ID>OUT_12</ID>1675 </output>
<output>
<ID>OUT_13</ID>1683 </output>
<output>
<ID>OUT_14</ID>1676 </output>
<output>
<ID>OUT_15</ID>1684 </output>
<output>
<ID>OUT_2</ID>1670 </output>
<output>
<ID>OUT_3</ID>1678 </output>
<output>
<ID>OUT_4</ID>1671 </output>
<output>
<ID>OUT_5</ID>1679 </output>
<output>
<ID>OUT_6</ID>1672 </output>
<output>
<ID>OUT_7</ID>1680 </output>
<output>
<ID>OUT_8</ID>1673 </output>
<output>
<ID>OUT_9</ID>1681 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1135</ID>
<type>AA_LABEL</type>
<position>568,1328</position>
<gparam>LABEL_TEXT 0 = ADD, 1 = AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1136</ID>
<type>AE_REGISTER8</type>
<position>450,1314</position>
<input>
<ID>IN_0</ID>1782 </input>
<input>
<ID>IN_1</ID>1781 </input>
<input>
<ID>IN_2</ID>1780 </input>
<input>
<ID>IN_3</ID>1779 </input>
<input>
<ID>IN_4</ID>1778 </input>
<input>
<ID>IN_5</ID>1777 </input>
<input>
<ID>IN_6</ID>1776 </input>
<input>
<ID>IN_7</ID>1775 </input>
<output>
<ID>OUT_0</ID>1746 </output>
<output>
<ID>OUT_1</ID>1745 </output>
<output>
<ID>OUT_2</ID>1744 </output>
<output>
<ID>OUT_3</ID>1743 </output>
<output>
<ID>OUT_4</ID>1742 </output>
<output>
<ID>OUT_5</ID>1741 </output>
<output>
<ID>OUT_6</ID>1740 </output>
<output>
<ID>OUT_7</ID>1739 </output>
<input>
<ID>clock</ID>1762 </input>
<input>
<ID>load</ID>1597 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1137</ID>
<type>AA_LABEL</type>
<position>612.5,1272.5</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1138</ID>
<type>AE_REGISTER8</type>
<position>450,1327</position>
<input>
<ID>IN_0</ID>1782 </input>
<input>
<ID>IN_1</ID>1781 </input>
<input>
<ID>IN_2</ID>1780 </input>
<input>
<ID>IN_3</ID>1779 </input>
<input>
<ID>IN_4</ID>1778 </input>
<input>
<ID>IN_5</ID>1777 </input>
<input>
<ID>IN_6</ID>1776 </input>
<input>
<ID>IN_7</ID>1775 </input>
<output>
<ID>OUT_0</ID>1761 </output>
<output>
<ID>OUT_1</ID>1752 </output>
<output>
<ID>OUT_2</ID>1751 </output>
<output>
<ID>OUT_3</ID>1586 </output>
<output>
<ID>OUT_4</ID>1750 </output>
<output>
<ID>OUT_5</ID>1749 </output>
<output>
<ID>OUT_6</ID>1748 </output>
<output>
<ID>OUT_7</ID>1747 </output>
<input>
<ID>clock</ID>1762 </input>
<input>
<ID>load</ID>1596 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1139</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1338</position>
<input>
<ID>IN_0</ID>1747 </input>
<input>
<ID>IN_1</ID>1739 </input>
<input>
<ID>IN_2</ID>1731 </input>
<input>
<ID>IN_3</ID>1785 </input>
<output>
<ID>OUT</ID>1753 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1140</ID>
<type>AA_LABEL</type>
<position>598.5,1301</position>
<gparam>LABEL_TEXT B0-B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1141</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1327</position>
<input>
<ID>IN_0</ID>1748 </input>
<input>
<ID>IN_1</ID>1740 </input>
<input>
<ID>IN_2</ID>1732 </input>
<input>
<ID>IN_3</ID>1725 </input>
<output>
<ID>OUT</ID>1754 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1142</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1316</position>
<input>
<ID>IN_0</ID>1749 </input>
<input>
<ID>IN_1</ID>1741 </input>
<input>
<ID>IN_2</ID>1733 </input>
<input>
<ID>IN_3</ID>1726 </input>
<output>
<ID>OUT</ID>1755 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1143</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1306.5</position>
<input>
<ID>IN_0</ID>1750 </input>
<input>
<ID>IN_1</ID>1742 </input>
<input>
<ID>IN_2</ID>1734 </input>
<input>
<ID>IN_3</ID>1727 </input>
<output>
<ID>OUT</ID>1756 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1144</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1295.5</position>
<input>
<ID>IN_0</ID>1586 </input>
<input>
<ID>IN_1</ID>1743 </input>
<input>
<ID>IN_2</ID>1735 </input>
<input>
<ID>IN_3</ID>1728 </input>
<output>
<ID>OUT</ID>1757 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1145</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1284.5</position>
<input>
<ID>IN_0</ID>1751 </input>
<input>
<ID>IN_1</ID>1744 </input>
<input>
<ID>IN_2</ID>1736 </input>
<input>
<ID>IN_3</ID>1556 </input>
<output>
<ID>OUT</ID>1758 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1146</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1274</position>
<input>
<ID>IN_0</ID>1752 </input>
<input>
<ID>IN_1</ID>1745 </input>
<input>
<ID>IN_2</ID>1737 </input>
<input>
<ID>IN_3</ID>1729 </input>
<output>
<ID>OUT</ID>1759 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1147</ID>
<type>AE_MUX_4x1</type>
<position>475.5,1263</position>
<input>
<ID>IN_0</ID>1761 </input>
<input>
<ID>IN_1</ID>1746 </input>
<input>
<ID>IN_2</ID>1738 </input>
<input>
<ID>IN_3</ID>1730 </input>
<output>
<ID>OUT</ID>1760 </output>
<input>
<ID>SEL_0</ID>1763 </input>
<input>
<ID>SEL_1</ID>1764 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1148</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>514,1304.5</position>
<input>
<ID>IN_0</ID>1760 </input>
<input>
<ID>IN_1</ID>1759 </input>
<input>
<ID>IN_2</ID>1758 </input>
<input>
<ID>IN_3</ID>1757 </input>
<input>
<ID>IN_4</ID>1756 </input>
<input>
<ID>IN_5</ID>1755 </input>
<input>
<ID>IN_6</ID>1754 </input>
<input>
<ID>IN_7</ID>1753 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1150</ID>
<type>AA_LABEL</type>
<position>598.5,1295</position>
<gparam>LABEL_TEXT A0-A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1151</ID>
<type>AA_LABEL</type>
<position>450,1334</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1152</ID>
<type>AA_LABEL</type>
<position>450,1321</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1153</ID>
<type>AA_LABEL</type>
<position>450,1307.5</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1154</ID>
<type>AA_LABEL</type>
<position>450,1294.5</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1157</ID>
<type>AE_MUX_4x1</type>
<position>488,1338</position>
<input>
<ID>IN_0</ID>1747 </input>
<input>
<ID>IN_1</ID>1739 </input>
<input>
<ID>IN_2</ID>1731 </input>
<input>
<ID>IN_3</ID>1785 </input>
<output>
<ID>OUT</ID>1765 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1158</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1318</position>
<input>
<ID>IN_0</ID>1708 </input>
<input>
<ID>IN_1</ID>1716 </input>
<output>
<ID>OUT</ID>1724 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1159</ID>
<type>AA_LABEL</type>
<position>598.5,1285</position>
<gparam>LABEL_TEXT B4-B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1160</ID>
<type>AE_MUX_4x1</type>
<position>488,1327</position>
<input>
<ID>IN_0</ID>1748 </input>
<input>
<ID>IN_1</ID>1740 </input>
<input>
<ID>IN_2</ID>1732 </input>
<input>
<ID>IN_3</ID>1725 </input>
<output>
<ID>OUT</ID>1766 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1161</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1313</position>
<input>
<ID>IN_0</ID>1707 </input>
<input>
<ID>IN_1</ID>1715 </input>
<output>
<ID>OUT</ID>1723 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1162</ID>
<type>AE_MUX_4x1</type>
<position>488,1316</position>
<input>
<ID>IN_0</ID>1749 </input>
<input>
<ID>IN_1</ID>1741 </input>
<input>
<ID>IN_2</ID>1733 </input>
<input>
<ID>IN_3</ID>1726 </input>
<output>
<ID>OUT</ID>1767 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1163</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1308</position>
<input>
<ID>IN_0</ID>1706 </input>
<input>
<ID>IN_1</ID>1714 </input>
<output>
<ID>OUT</ID>1722 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1164</ID>
<type>AE_MUX_4x1</type>
<position>488,1306.5</position>
<input>
<ID>IN_0</ID>1750 </input>
<input>
<ID>IN_1</ID>1742 </input>
<input>
<ID>IN_2</ID>1734 </input>
<input>
<ID>IN_3</ID>1727 </input>
<output>
<ID>OUT</ID>1768 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1165</ID>
<type>AE_MUX_4x1</type>
<position>488,1295.5</position>
<input>
<ID>IN_0</ID>1586 </input>
<input>
<ID>IN_1</ID>1743 </input>
<input>
<ID>IN_2</ID>1735 </input>
<input>
<ID>IN_3</ID>1728 </input>
<output>
<ID>OUT</ID>1769 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1166</ID>
<type>AE_MUX_4x1</type>
<position>488,1284.5</position>
<input>
<ID>IN_0</ID>1751 </input>
<input>
<ID>IN_1</ID>1744 </input>
<input>
<ID>IN_2</ID>1736 </input>
<input>
<ID>IN_3</ID>1556 </input>
<output>
<ID>OUT</ID>1770 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1167</ID>
<type>AE_MUX_4x1</type>
<position>488,1274</position>
<input>
<ID>IN_0</ID>1752 </input>
<input>
<ID>IN_1</ID>1745 </input>
<input>
<ID>IN_2</ID>1737 </input>
<input>
<ID>IN_3</ID>1729 </input>
<output>
<ID>OUT</ID>1771 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1168</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1303</position>
<input>
<ID>IN_0</ID>1705 </input>
<input>
<ID>IN_1</ID>1713 </input>
<output>
<ID>OUT</ID>1721 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1169</ID>
<type>AA_LABEL</type>
<position>599.5,1278</position>
<gparam>LABEL_TEXT A4-A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1170</ID>
<type>AE_MUX_4x1</type>
<position>488,1263</position>
<input>
<ID>IN_0</ID>1761 </input>
<input>
<ID>IN_1</ID>1746 </input>
<input>
<ID>IN_2</ID>1738 </input>
<input>
<ID>IN_3</ID>1730 </input>
<output>
<ID>OUT</ID>1772 </output>
<input>
<ID>SEL_0</ID>1773 </input>
<input>
<ID>SEL_1</ID>1774 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1171</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1298</position>
<input>
<ID>IN_0</ID>1704 </input>
<input>
<ID>IN_1</ID>1712 </input>
<output>
<ID>OUT</ID>1720 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1172</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>514,1294.5</position>
<input>
<ID>IN_0</ID>1772 </input>
<input>
<ID>IN_1</ID>1771 </input>
<input>
<ID>IN_2</ID>1770 </input>
<input>
<ID>IN_3</ID>1769 </input>
<input>
<ID>IN_4</ID>1768 </input>
<input>
<ID>IN_5</ID>1767 </input>
<input>
<ID>IN_6</ID>1766 </input>
<input>
<ID>IN_7</ID>1765 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 52</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1173</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1293</position>
<input>
<ID>IN_0</ID>1703 </input>
<input>
<ID>IN_1</ID>1711 </input>
<output>
<ID>OUT</ID>1719 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1174</ID>
<type>DE_TO</type>
<position>756,1318.5</position>
<input>
<ID>IN_0</ID>1515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BR</lparam></gate>
<gate>
<ID>1176</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1288</position>
<input>
<ID>IN_0</ID>1702 </input>
<input>
<ID>IN_1</ID>1710 </input>
<output>
<ID>OUT</ID>1718 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1177</ID>
<type>AE_FULLADDER_4BIT</type>
<position>702.5,1350</position>
<input>
<ID>IN_0</ID>1532 </input>
<input>
<ID>IN_1</ID>1534 </input>
<input>
<ID>IN_2</ID>1536 </input>
<input>
<ID>IN_3</ID>1553 </input>
<input>
<ID>IN_B_0</ID>1998 </input>
<output>
<ID>OUT_0</ID>1615 </output>
<output>
<ID>OUT_1</ID>1620 </output>
<output>
<ID>OUT_2</ID>1621 </output>
<output>
<ID>OUT_3</ID>1622 </output>
<output>
<ID>carry_out</ID>1516 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1178</ID>
<type>AA_MUX_2x1</type>
<position>630.5,1283</position>
<input>
<ID>IN_0</ID>1701 </input>
<input>
<ID>IN_1</ID>1709 </input>
<output>
<ID>OUT</ID>1717 </output>
<input>
<ID>SEL_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1179</ID>
<type>AE_FULLADDER_4BIT</type>
<position>702.5,1334</position>
<input>
<ID>IN_0</ID>1602 </input>
<input>
<ID>IN_1</ID>1603 </input>
<input>
<ID>IN_2</ID>1608 </input>
<input>
<ID>IN_3</ID>1609 </input>
<output>
<ID>OUT_0</ID>1664 </output>
<output>
<ID>OUT_1</ID>1783 </output>
<output>
<ID>OUT_2</ID>1837 </output>
<output>
<ID>OUT_3</ID>1997 </output>
<input>
<ID>carry_in</ID>1516 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1180</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>676.5,1299.5</position>
<input>
<ID>IN_0</ID>1717 </input>
<input>
<ID>IN_1</ID>1718 </input>
<input>
<ID>IN_2</ID>1719 </input>
<input>
<ID>IN_3</ID>1720 </input>
<input>
<ID>IN_4</ID>1721 </input>
<input>
<ID>IN_5</ID>1722 </input>
<input>
<ID>IN_6</ID>1723 </input>
<input>
<ID>IN_7</ID>1724 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 104</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1181</ID>
<type>BA_DECODER_2x4</type>
<position>435,1342.5</position>
<input>
<ID>ENABLE</ID>1044 </input>
<input>
<ID>IN_0</ID>1601 </input>
<input>
<ID>IN_1</ID>1600 </input>
<output>
<ID>OUT_0</ID>1596 </output>
<output>
<ID>OUT_1</ID>1597 </output>
<output>
<ID>OUT_2</ID>1598 </output>
<output>
<ID>OUT_3</ID>1599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1182</ID>
<type>AA_LABEL</type>
<position>633,1280</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1184</ID>
<type>AA_LABEL</type>
<position>633,1322</position>
<gparam>LABEL_TEXT A7/B7</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1185</ID>
<type>AA_AND2</type>
<position>600.5,1305</position>
<input>
<ID>IN_0</ID>1686 </input>
<input>
<ID>IN_1</ID>1685 </input>
<output>
<ID>OUT</ID>1709 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1187</ID>
<type>GA_LED</type>
<position>644.5,1291</position>
<input>
<ID>N_in2</ID>1724 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1189</ID>
<type>GA_LED</type>
<position>647,1291</position>
<input>
<ID>N_in2</ID>1723 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1191</ID>
<type>GA_LED</type>
<position>649.5,1291</position>
<input>
<ID>N_in2</ID>1722 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1192</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>532,1313.5</position>
<input>
<ID>ENABLE_0</ID>1519 </input>
<input>
<ID>IN_0</ID>1760 </input>
<input>
<ID>IN_1</ID>1759 </input>
<input>
<ID>IN_2</ID>1758 </input>
<input>
<ID>IN_3</ID>1757 </input>
<input>
<ID>IN_4</ID>1756 </input>
<input>
<ID>IN_5</ID>1755 </input>
<input>
<ID>IN_6</ID>1754 </input>
<input>
<ID>IN_7</ID>1753 </input>
<output>
<ID>OUT_0</ID>1790 </output>
<output>
<ID>OUT_1</ID>1789 </output>
<output>
<ID>OUT_2</ID>1788 </output>
<output>
<ID>OUT_3</ID>2082 </output>
<output>
<ID>OUT_4</ID>2083 </output>
<output>
<ID>OUT_5</ID>2084 </output>
<output>
<ID>OUT_6</ID>2085 </output>
<output>
<ID>OUT_7</ID>2089 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1193</ID>
<type>GA_LED</type>
<position>652,1291</position>
<input>
<ID>N_in2</ID>1721 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1194</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>532,1286.5</position>
<input>
<ID>ENABLE_0</ID>1784 </input>
<input>
<ID>IN_0</ID>1772 </input>
<input>
<ID>IN_1</ID>1771 </input>
<input>
<ID>IN_2</ID>1770 </input>
<input>
<ID>IN_3</ID>1769 </input>
<input>
<ID>IN_4</ID>1768 </input>
<input>
<ID>IN_5</ID>1767 </input>
<input>
<ID>IN_6</ID>1766 </input>
<input>
<ID>IN_7</ID>1765 </input>
<output>
<ID>OUT_0</ID>1798 </output>
<output>
<ID>OUT_1</ID>1797 </output>
<output>
<ID>OUT_2</ID>1796 </output>
<output>
<ID>OUT_3</ID>1795 </output>
<output>
<ID>OUT_4</ID>1794 </output>
<output>
<ID>OUT_5</ID>1793 </output>
<output>
<ID>OUT_6</ID>1792 </output>
<output>
<ID>OUT_7</ID>1791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1195</ID>
<type>GA_LED</type>
<position>654.5,1291</position>
<input>
<ID>N_in2</ID>1720 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1196</ID>
<type>AA_AND2</type>
<position>605.5,1308.5</position>
<input>
<ID>IN_0</ID>1688 </input>
<input>
<ID>IN_1</ID>1687 </input>
<output>
<ID>OUT</ID>1710 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1197</ID>
<type>AA_LABEL</type>
<position>532,1308.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1198</ID>
<type>GA_LED</type>
<position>657,1291</position>
<input>
<ID>N_in2</ID>1719 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1199</ID>
<type>AA_LABEL</type>
<position>505.5,1301</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1200</ID>
<type>GA_LED</type>
<position>659.5,1291</position>
<input>
<ID>N_in2</ID>1718 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1201</ID>
<type>AA_LABEL</type>
<position>532,1281.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1202</ID>
<type>GA_LED</type>
<position>662,1291</position>
<input>
<ID>N_in2</ID>1717 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam></gate>
<gate>
<ID>1203</ID>
<type>AA_LABEL</type>
<position>505.5,1299.5</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1204</ID>
<type>AA_LABEL</type>
<position>662,1289</position>
<gparam>LABEL_TEXT F0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1205</ID>
<type>EE_VDD</type>
<position>532,1293.5</position>
<output>
<ID>OUT_0</ID>1784 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1206</ID>
<type>AA_LABEL</type>
<position>659.5,1289</position>
<gparam>LABEL_TEXT F1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1207</ID>
<type>BA_DECODER_2x4</type>
<position>579,1330</position>
<input>
<ID>ENABLE</ID>2023 </input>
<input>
<ID>IN_0</ID>1665 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<output>
<ID>OUT_1</ID>1667 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1208</ID>
<type>AA_LABEL</type>
<position>657,1289</position>
<gparam>LABEL_TEXT F2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1210</ID>
<type>AA_LABEL</type>
<position>654.5,1289</position>
<gparam>LABEL_TEXT F3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1211</ID>
<type>AA_AND2</type>
<position>600.5,1312</position>
<input>
<ID>IN_0</ID>1690 </input>
<input>
<ID>IN_1</ID>1689 </input>
<output>
<ID>OUT</ID>1711 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1213</ID>
<type>AA_LABEL</type>
<position>652,1289</position>
<gparam>LABEL_TEXT F4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1215</ID>
<type>AE_FULLADDER_4BIT</type>
<position>605,1295</position>
<input>
<ID>IN_0</ID>1677 </input>
<input>
<ID>IN_1</ID>1678 </input>
<input>
<ID>IN_2</ID>1679 </input>
<input>
<ID>IN_3</ID>1680 </input>
<input>
<ID>IN_B_0</ID>1669 </input>
<input>
<ID>IN_B_1</ID>1670 </input>
<input>
<ID>IN_B_2</ID>1671 </input>
<input>
<ID>IN_B_3</ID>1672 </input>
<output>
<ID>OUT_0</ID>1701 </output>
<output>
<ID>OUT_1</ID>1702 </output>
<output>
<ID>OUT_2</ID>1703 </output>
<output>
<ID>OUT_3</ID>1704 </output>
<output>
<ID>carry_out</ID>1668 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1216</ID>
<type>AE_FULLADDER_4BIT</type>
<position>605,1278.5</position>
<input>
<ID>IN_0</ID>1681 </input>
<input>
<ID>IN_1</ID>1682 </input>
<input>
<ID>IN_2</ID>1683 </input>
<input>
<ID>IN_3</ID>1684 </input>
<input>
<ID>IN_B_0</ID>1673 </input>
<input>
<ID>IN_B_1</ID>1674 </input>
<input>
<ID>IN_B_2</ID>1675 </input>
<input>
<ID>IN_B_3</ID>1676 </input>
<output>
<ID>OUT_0</ID>1705 </output>
<output>
<ID>OUT_1</ID>1706 </output>
<output>
<ID>OUT_2</ID>1707 </output>
<output>
<ID>OUT_3</ID>1708 </output>
<input>
<ID>carry_in</ID>1668 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1217</ID>
<type>AA_LABEL</type>
<position>649.5,1289</position>
<gparam>LABEL_TEXT F5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1218</ID>
<type>AA_LABEL</type>
<position>612.5,1301.5</position>
<gparam>LABEL_TEXT A0/B0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1219</ID>
<type>AA_LABEL</type>
<position>647,1289</position>
<gparam>LABEL_TEXT F6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1220</ID>
<type>DE_TO</type>
<position>559,1405.5</position>
<input>
<ID>IN_0</ID>1831 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC7</lparam></gate>
<gate>
<ID>1221</ID>
<type>DE_TO</type>
<position>559,1403.5</position>
<input>
<ID>IN_0</ID>1832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC6</lparam></gate>
<gate>
<ID>1222</ID>
<type>AA_LABEL</type>
<position>644.5,1289</position>
<gparam>LABEL_TEXT F7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1223</ID>
<type>DE_TO</type>
<position>559,1401.5</position>
<input>
<ID>IN_0</ID>1833 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC5</lparam></gate>
<gate>
<ID>1225</ID>
<type>AA_AND2</type>
<position>605.5,1315.5</position>
<input>
<ID>IN_0</ID>1692 </input>
<input>
<ID>IN_1</ID>1691 </input>
<output>
<ID>OUT</ID>1712 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1226</ID>
<type>DE_TO</type>
<position>559,1399.5</position>
<input>
<ID>IN_0</ID>1834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC4</lparam></gate>
<gate>
<ID>1228</ID>
<type>DE_TO</type>
<position>559,1397.5</position>
<input>
<ID>IN_0</ID>1835 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC3</lparam></gate>
<gate>
<ID>1229</ID>
<type>AA_LABEL</type>
<position>574,1334</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1230</ID>
<type>DE_TO</type>
<position>559,1395.5</position>
<input>
<ID>IN_0</ID>1836 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC2</lparam></gate>
<gate>
<ID>1232</ID>
<type>DE_TO</type>
<position>559,1393.5</position>
<input>
<ID>IN_0</ID>1968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC1</lparam></gate>
<gate>
<ID>1233</ID>
<type>DE_TO</type>
<position>559,1391.5</position>
<input>
<ID>IN_0</ID>1838 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC0</lparam></gate>
<gate>
<ID>1234</ID>
<type>AA_AND2</type>
<position>600.5,1319</position>
<input>
<ID>IN_0</ID>1694 </input>
<input>
<ID>IN_1</ID>1693 </input>
<output>
<ID>OUT</ID>1713 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1235</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>430,1362</position>
<input>
<ID>ENABLE_0</ID>2090 </input>
<input>
<ID>IN_0</ID>1845 </input>
<input>
<ID>IN_1</ID>1844 </input>
<input>
<ID>IN_2</ID>2078 </input>
<input>
<ID>IN_3</ID>2079 </input>
<input>
<ID>IN_4</ID>1841 </input>
<input>
<ID>IN_5</ID>1856 </input>
<input>
<ID>IN_6</ID>1840 </input>
<input>
<ID>IN_7</ID>1839 </input>
<output>
<ID>OUT_0</ID>1855 </output>
<output>
<ID>OUT_1</ID>1854 </output>
<output>
<ID>OUT_2</ID>1853 </output>
<output>
<ID>OUT_3</ID>1852 </output>
<output>
<ID>OUT_4</ID>1851 </output>
<output>
<ID>OUT_5</ID>1850 </output>
<output>
<ID>OUT_6</ID>1849 </output>
<output>
<ID>OUT_7</ID>1848 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1236</ID>
<type>DA_FROM</type>
<position>419,1365.5</position>
<input>
<ID>IN_0</ID>1839 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC7</lparam></gate>
<gate>
<ID>1237</ID>
<type>DA_FROM</type>
<position>419,1363.5</position>
<input>
<ID>IN_0</ID>1840 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC6</lparam></gate>
<gate>
<ID>1238</ID>
<type>DA_FROM</type>
<position>419,1361.5</position>
<input>
<ID>IN_0</ID>1856 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC5</lparam></gate>
<gate>
<ID>1239</ID>
<type>DA_FROM</type>
<position>419,1359.5</position>
<input>
<ID>IN_0</ID>1841 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC4</lparam></gate>
<gate>
<ID>1240</ID>
<type>DA_FROM</type>
<position>419,1355.5</position>
<input>
<ID>IN_0</ID>2078 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC2</lparam></gate>
<gate>
<ID>1241</ID>
<type>DA_FROM</type>
<position>419,1357.5</position>
<input>
<ID>IN_0</ID>2079 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC3</lparam></gate>
<gate>
<ID>1242</ID>
<type>DA_FROM</type>
<position>419,1353.5</position>
<input>
<ID>IN_0</ID>1844 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC1</lparam></gate>
<gate>
<ID>1243</ID>
<type>DA_FROM</type>
<position>419,1351.5</position>
<input>
<ID>IN_0</ID>1845 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC0</lparam></gate>
<gate>
<ID>1244</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>447,1362.5</position>
<input>
<ID>ENABLE_0</ID>1895 </input>
<input>
<ID>IN_0</ID>1855 </input>
<input>
<ID>IN_1</ID>1854 </input>
<input>
<ID>IN_2</ID>1853 </input>
<input>
<ID>IN_3</ID>1852 </input>
<input>
<ID>IN_4</ID>1851 </input>
<input>
<ID>IN_5</ID>1850 </input>
<input>
<ID>IN_6</ID>1849 </input>
<input>
<ID>IN_7</ID>1848 </input>
<output>
<ID>OUT_0</ID>1865 </output>
<output>
<ID>OUT_1</ID>1864 </output>
<output>
<ID>OUT_2</ID>1863 </output>
<output>
<ID>OUT_3</ID>1862 </output>
<output>
<ID>OUT_4</ID>1861 </output>
<output>
<ID>OUT_5</ID>1860 </output>
<output>
<ID>OUT_6</ID>1859 </output>
<output>
<ID>OUT_7</ID>1858 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1246</ID>
<type>DA_FROM</type>
<position>696,1327.5</position>
<input>
<ID>IN_0</ID>1609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC7</lparam></gate>
<gate>
<ID>1247</ID>
<type>DE_TO</type>
<position>457,1373</position>
<input>
<ID>IN_0</ID>1858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR7</lparam></gate>
<gate>
<ID>1248</ID>
<type>EE_VDD</type>
<position>447,1369.5</position>
<output>
<ID>OUT_0</ID>1895 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1249</ID>
<type>DE_TO</type>
<position>457,1371</position>
<input>
<ID>IN_0</ID>1859 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR6</lparam></gate>
<gate>
<ID>1250</ID>
<type>DE_TO</type>
<position>457,1369</position>
<input>
<ID>IN_0</ID>1860 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR5</lparam></gate>
<gate>
<ID>1251</ID>
<type>DE_TO</type>
<position>457,1367</position>
<input>
<ID>IN_0</ID>1861 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR4</lparam></gate>
<gate>
<ID>1252</ID>
<type>DE_TO</type>
<position>457,1365</position>
<input>
<ID>IN_0</ID>1862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR3</lparam></gate>
<gate>
<ID>1253</ID>
<type>DE_TO</type>
<position>457,1363</position>
<input>
<ID>IN_0</ID>1863 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR2</lparam></gate>
<gate>
<ID>1254</ID>
<type>DE_TO</type>
<position>457,1361</position>
<input>
<ID>IN_0</ID>1864 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR1</lparam></gate>
<gate>
<ID>1255</ID>
<type>DE_TO</type>
<position>457,1359</position>
<input>
<ID>IN_0</ID>1865 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR0</lparam></gate>
<gate>
<ID>1256</ID>
<type>DA_FROM</type>
<position>560.5,1382.5</position>
<input>
<ID>IN_0</ID>1866 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR7</lparam></gate>
<gate>
<ID>1257</ID>
<type>DA_FROM</type>
<position>560.5,1380.5</position>
<input>
<ID>IN_0</ID>1867 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR6</lparam></gate>
<gate>
<ID>1259</ID>
<type>AA_LABEL</type>
<position>573.5,1397.5</position>
<gparam>LABEL_TEXT MAR Load Control</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1260</ID>
<type>DA_FROM</type>
<position>560.5,1374.5</position>
<input>
<ID>IN_0</ID>1871 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR3</lparam></gate>
<gate>
<ID>1261</ID>
<type>DA_FROM</type>
<position>560.5,1378.5</position>
<input>
<ID>IN_0</ID>1873 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR5</lparam></gate>
<gate>
<ID>1262</ID>
<type>DA_FROM</type>
<position>560.5,1372.5</position>
<input>
<ID>IN_0</ID>1870 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR2</lparam></gate>
<gate>
<ID>1263</ID>
<type>DA_FROM</type>
<position>560.5,1370.5</position>
<input>
<ID>IN_0</ID>1869 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR1</lparam></gate>
<gate>
<ID>1264</ID>
<type>DA_FROM</type>
<position>560.5,1368.5</position>
<input>
<ID>IN_0</ID>1868 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR0</lparam></gate>
<gate>
<ID>1265</ID>
<type>DA_FROM</type>
<position>560.5,1376.5</position>
<input>
<ID>IN_0</ID>1872 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR4</lparam></gate>
<gate>
<ID>1266</ID>
<type>AA_TOGGLE</type>
<position>567.5,1395.5</position>
<output>
<ID>OUT_0</ID>1874 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1267</ID>
<type>DA_FROM</type>
<position>696,1329.5</position>
<input>
<ID>IN_0</ID>1608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC6</lparam></gate>
<gate>
<ID>1268</ID>
<type>AE_FULLADDER_4BIT</type>
<position>698.5,1386</position>
<input>
<ID>IN_0</ID>1886 </input>
<input>
<ID>IN_1</ID>1887 </input>
<input>
<ID>IN_2</ID>1888 </input>
<input>
<ID>IN_3</ID>1889 </input>
<input>
<ID>IN_B_0</ID>1882 </input>
<input>
<ID>IN_B_1</ID>1883 </input>
<input>
<ID>IN_B_2</ID>1884 </input>
<input>
<ID>IN_B_3</ID>1885 </input>
<output>
<ID>OUT_0</ID>1896 </output>
<output>
<ID>OUT_1</ID>1897 </output>
<output>
<ID>OUT_2</ID>1898 </output>
<output>
<ID>OUT_3</ID>1899 </output>
<output>
<ID>carry_out</ID>1876 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1269</ID>
<type>AE_FULLADDER_4BIT</type>
<position>698.5,1370</position>
<input>
<ID>IN_0</ID>1890 </input>
<input>
<ID>IN_1</ID>1891 </input>
<input>
<ID>IN_2</ID>1892 </input>
<input>
<ID>IN_3</ID>1893 </input>
<input>
<ID>IN_B_0</ID>1881 </input>
<input>
<ID>IN_B_1</ID>1880 </input>
<input>
<ID>IN_B_2</ID>1879 </input>
<input>
<ID>IN_B_3</ID>1878 </input>
<output>
<ID>OUT_0</ID>1900 </output>
<output>
<ID>OUT_1</ID>1901 </output>
<output>
<ID>OUT_2</ID>1902 </output>
<output>
<ID>OUT_3</ID>1903 </output>
<input>
<ID>carry_in</ID>1876 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1270</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>636,1375</position>
<input>
<ID>ENABLE_0</ID>1943 </input>
<input>
<ID>IN_0</ID>1616 </input>
<input>
<ID>IN_1</ID>1614 </input>
<input>
<ID>IN_2</ID>1613 </input>
<input>
<ID>IN_3</ID>1612 </input>
<output>
<ID>OUT_0</ID>1882 </output>
<output>
<ID>OUT_1</ID>1883 </output>
<output>
<ID>OUT_2</ID>1884 </output>
<output>
<ID>OUT_3</ID>1877 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1271</ID>
<type>DE_TO</type>
<position>642.5,1374.5</position>
<input>
<ID>IN_0</ID>1877 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1272</ID>
<type>DA_FROM</type>
<position>691.5,1372</position>
<input>
<ID>IN_0</ID>1878 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1273</ID>
<type>DA_FROM</type>
<position>691.5,1374</position>
<input>
<ID>IN_0</ID>1879 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1274</ID>
<type>DA_FROM</type>
<position>691.5,1376</position>
<input>
<ID>IN_0</ID>1880 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1275</ID>
<type>DA_FROM</type>
<position>691.5,1378</position>
<input>
<ID>IN_0</ID>1881 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1276</ID>
<type>DA_FROM</type>
<position>691.5,1388</position>
<input>
<ID>IN_0</ID>1885 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID signbit</lparam></gate>
<gate>
<ID>1277</ID>
<type>DA_FROM</type>
<position>691.5,1364</position>
<input>
<ID>IN_0</ID>1893 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC7</lparam></gate>
<gate>
<ID>1278</ID>
<type>DA_FROM</type>
<position>691.5,1366</position>
<input>
<ID>IN_0</ID>1892 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC6</lparam></gate>
<gate>
<ID>1279</ID>
<type>DA_FROM</type>
<position>691.5,1368</position>
<input>
<ID>IN_0</ID>1891 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC5</lparam></gate>
<gate>
<ID>1280</ID>
<type>DA_FROM</type>
<position>691.5,1370</position>
<input>
<ID>IN_0</ID>1890 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC4</lparam></gate>
<gate>
<ID>1281</ID>
<type>DA_FROM</type>
<position>691.5,1382</position>
<input>
<ID>IN_0</ID>1888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC2</lparam></gate>
<gate>
<ID>1282</ID>
<type>DA_FROM</type>
<position>691.5,1380</position>
<input>
<ID>IN_0</ID>1889 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC3</lparam></gate>
<gate>
<ID>1283</ID>
<type>DA_FROM</type>
<position>691.5,1384</position>
<input>
<ID>IN_0</ID>1887 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC1</lparam></gate>
<gate>
<ID>1284</ID>
<type>DA_FROM</type>
<position>691.5,1386</position>
<input>
<ID>IN_0</ID>1886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC0</lparam></gate>
<gate>
<ID>1285</ID>
<type>DA_FROM</type>
<position>696,1331.5</position>
<input>
<ID>IN_0</ID>1603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC5</lparam></gate>
<gate>
<ID>1286</ID>
<type>AA_INVERTER</type>
<position>597,1382.5</position>
<input>
<ID>IN_0</ID>1645 </input>
<output>
<ID>OUT_0</ID>1786 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1288</ID>
<type>DA_FROM</type>
<position>696,1333.5</position>
<input>
<ID>IN_0</ID>1602 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC4</lparam></gate>
<gate>
<ID>1289</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>572.5,1313.5</position>
<input>
<ID>ENABLE_0</ID>1618 </input>
<input>
<ID>IN_0</ID>1798 </input>
<input>
<ID>IN_1</ID>1790 </input>
<input>
<ID>IN_10</ID>1793 </input>
<input>
<ID>IN_11</ID>2084 </input>
<input>
<ID>IN_12</ID>1792 </input>
<input>
<ID>IN_13</ID>2085 </input>
<input>
<ID>IN_14</ID>1791 </input>
<input>
<ID>IN_15</ID>2089 </input>
<input>
<ID>IN_2</ID>1797 </input>
<input>
<ID>IN_3</ID>1789 </input>
<input>
<ID>IN_4</ID>1796 </input>
<input>
<ID>IN_5</ID>1788 </input>
<input>
<ID>IN_6</ID>1795 </input>
<input>
<ID>IN_7</ID>2082 </input>
<input>
<ID>IN_8</ID>1794 </input>
<input>
<ID>IN_9</ID>2083 </input>
<output>
<ID>OUT_0</ID>1822 </output>
<output>
<ID>OUT_1</ID>1815 </output>
<output>
<ID>OUT_10</ID>1827 </output>
<output>
<ID>OUT_11</ID>1828 </output>
<output>
<ID>OUT_12</ID>1825 </output>
<output>
<ID>OUT_13</ID>1823 </output>
<output>
<ID>OUT_14</ID>1826 </output>
<output>
<ID>OUT_15</ID>1830 </output>
<output>
<ID>OUT_2</ID>1819 </output>
<output>
<ID>OUT_3</ID>1818 </output>
<output>
<ID>OUT_4</ID>1816 </output>
<output>
<ID>OUT_5</ID>1817 </output>
<output>
<ID>OUT_6</ID>1820 </output>
<output>
<ID>OUT_7</ID>1821 </output>
<output>
<ID>OUT_8</ID>1829 </output>
<output>
<ID>OUT_9</ID>1824 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1290</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>572.5,1290.5</position>
<input>
<ID>ENABLE_0</ID>1617 </input>
<input>
<ID>IN_0</ID>1798 </input>
<input>
<ID>IN_1</ID>1790 </input>
<input>
<ID>IN_10</ID>1793 </input>
<input>
<ID>IN_11</ID>2084 </input>
<input>
<ID>IN_12</ID>1792 </input>
<input>
<ID>IN_13</ID>2085 </input>
<input>
<ID>IN_14</ID>1791 </input>
<input>
<ID>IN_15</ID>2089 </input>
<input>
<ID>IN_2</ID>1797 </input>
<input>
<ID>IN_3</ID>1789 </input>
<input>
<ID>IN_4</ID>1796 </input>
<input>
<ID>IN_5</ID>1788 </input>
<input>
<ID>IN_6</ID>1795 </input>
<input>
<ID>IN_7</ID>2082 </input>
<input>
<ID>IN_8</ID>1794 </input>
<input>
<ID>IN_9</ID>2083 </input>
<output>
<ID>OUT_0</ID>1799 </output>
<output>
<ID>OUT_1</ID>1801 </output>
<output>
<ID>OUT_10</ID>1808 </output>
<output>
<ID>OUT_11</ID>1810 </output>
<output>
<ID>OUT_12</ID>1811 </output>
<output>
<ID>OUT_13</ID>1813 </output>
<output>
<ID>OUT_14</ID>1812 </output>
<output>
<ID>OUT_15</ID>1814 </output>
<output>
<ID>OUT_2</ID>1800 </output>
<output>
<ID>OUT_3</ID>1802 </output>
<output>
<ID>OUT_4</ID>1803 </output>
<output>
<ID>OUT_5</ID>1804 </output>
<output>
<ID>OUT_6</ID>1806 </output>
<output>
<ID>OUT_7</ID>1805 </output>
<output>
<ID>OUT_8</ID>1809 </output>
<output>
<ID>OUT_9</ID>1807 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1292</ID>
<type>DA_FROM</type>
<position>696,1345.5</position>
<input>
<ID>IN_0</ID>1536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC2</lparam></gate>
<gate>
<ID>1295</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>404,1329</position>
<input>
<ID>ENABLE_0</ID>2001 </input>
<input>
<ID>IN_0</ID>2094 </input>
<output>
<ID>OUT_0</ID>1763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1296</ID>
<type>AA_AND2</type>
<position>656,1344</position>
<input>
<ID>IN_0</ID>1605 </input>
<input>
<ID>IN_1</ID>1606 </input>
<output>
<ID>OUT</ID>1029 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1297</ID>
<type>DA_FROM</type>
<position>696,1343.5</position>
<input>
<ID>IN_0</ID>1553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC3</lparam></gate>
<gate>
<ID>1298</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>427,1309.5</position>
<input>
<ID>ENABLE_0</ID>1996 </input>
<input>
<ID>IN_0</ID>2095 </input>
<output>
<ID>OUT_0</ID>1601 </output>
<output>
<ID>OUT_1</ID>1600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1299</ID>
<type>DA_FROM</type>
<position>696,1347.5</position>
<input>
<ID>IN_0</ID>1534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC1</lparam></gate>
<gate>
<ID>1300</ID>
<type>DA_FROM</type>
<position>696,1349.5</position>
<input>
<ID>IN_0</ID>1532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC0</lparam></gate>
<gate>
<ID>1302</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>430,1377.5</position>
<input>
<ID>ENABLE_0</ID>1963 </input>
<input>
<ID>IN_0</ID>1911 </input>
<input>
<ID>IN_1</ID>1910 </input>
<input>
<ID>IN_2</ID>1909 </input>
<input>
<ID>IN_3</ID>1908 </input>
<input>
<ID>IN_4</ID>1907 </input>
<input>
<ID>IN_5</ID>1906 </input>
<input>
<ID>IN_6</ID>1905 </input>
<input>
<ID>IN_7</ID>1904 </input>
<output>
<ID>OUT_0</ID>1855 </output>
<output>
<ID>OUT_1</ID>1854 </output>
<output>
<ID>OUT_2</ID>1853 </output>
<output>
<ID>OUT_3</ID>1852 </output>
<output>
<ID>OUT_4</ID>1851 </output>
<output>
<ID>OUT_5</ID>1850 </output>
<output>
<ID>OUT_6</ID>1849 </output>
<output>
<ID>OUT_7</ID>1848 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1303</ID>
<type>AA_LABEL</type>
<position>701.5,1360</position>
<gparam>LABEL_TEXT PC + 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1304</ID>
<type>AA_LABEL</type>
<position>698,1397</position>
<gparam>LABEL_TEXT PC + off4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1306</ID>
<type>DE_TO</type>
<position>705,1389</position>
<input>
<ID>IN_0</ID>1896 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-0</lparam></gate>
<gate>
<ID>1307</ID>
<type>DE_TO</type>
<position>705,1387</position>
<input>
<ID>IN_0</ID>1897 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-1</lparam></gate>
<gate>
<ID>1308</ID>
<type>DE_TO</type>
<position>705,1385</position>
<input>
<ID>IN_0</ID>1898 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-2</lparam></gate>
<gate>
<ID>1309</ID>
<type>DE_TO</type>
<position>705,1383</position>
<input>
<ID>IN_0</ID>1899 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-3</lparam></gate>
<gate>
<ID>1310</ID>
<type>DE_TO</type>
<position>705,1373</position>
<input>
<ID>IN_0</ID>1900 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-4</lparam></gate>
<gate>
<ID>1311</ID>
<type>DE_TO</type>
<position>705,1371</position>
<input>
<ID>IN_0</ID>1901 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-5</lparam></gate>
<gate>
<ID>1312</ID>
<type>DE_TO</type>
<position>705,1369</position>
<input>
<ID>IN_0</ID>1902 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-6</lparam></gate>
<gate>
<ID>1313</ID>
<type>DE_TO</type>
<position>705,1367</position>
<input>
<ID>IN_0</ID>1903 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-7</lparam></gate>
<gate>
<ID>1314</ID>
<type>DE_TO</type>
<position>709,1353</position>
<input>
<ID>IN_0</ID>1615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-0</lparam></gate>
<gate>
<ID>1316</ID>
<type>DE_TO</type>
<position>709,1351</position>
<input>
<ID>IN_0</ID>1620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-1</lparam></gate>
<gate>
<ID>1317</ID>
<type>DA_FROM</type>
<position>421,1388</position>
<input>
<ID>IN_0</ID>1904 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-7</lparam></gate>
<gate>
<ID>1319</ID>
<type>DA_FROM</type>
<position>421,1386</position>
<input>
<ID>IN_0</ID>1905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-6</lparam></gate>
<gate>
<ID>1320</ID>
<type>DA_FROM</type>
<position>421,1384</position>
<input>
<ID>IN_0</ID>1906 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-5</lparam></gate>
<gate>
<ID>1321</ID>
<type>DA_FROM</type>
<position>421,1382</position>
<input>
<ID>IN_0</ID>1907 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-4</lparam></gate>
<gate>
<ID>1322</ID>
<type>DA_FROM</type>
<position>421,1380</position>
<input>
<ID>IN_0</ID>1908 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-3</lparam></gate>
<gate>
<ID>1323</ID>
<type>DA_FROM</type>
<position>421,1378</position>
<input>
<ID>IN_0</ID>1909 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-2</lparam></gate>
<gate>
<ID>1324</ID>
<type>DA_FROM</type>
<position>421,1376</position>
<input>
<ID>IN_0</ID>1910 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-1</lparam></gate>
<gate>
<ID>1325</ID>
<type>DA_FROM</type>
<position>421,1374</position>
<input>
<ID>IN_0</ID>1911 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff4-0</lparam></gate>
<gate>
<ID>1326</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>636.5,1392</position>
<input>
<ID>ENABLE_0</ID>1944 </input>
<input>
<ID>IN_0</ID>1616 </input>
<input>
<ID>IN_1</ID>1614 </input>
<input>
<ID>IN_2</ID>1613 </input>
<output>
<ID>OUT_0</ID>1941 </output>
<output>
<ID>OUT_1</ID>1942 </output>
<output>
<ID>OUT_2</ID>1940 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1327</ID>
<type>DE_TO</type>
<position>709,1349</position>
<input>
<ID>IN_0</ID>1621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-2</lparam></gate>
<gate>
<ID>1328</ID>
<type>AE_FULLADDER_4BIT</type>
<position>668.5,1412</position>
<input>
<ID>IN_0</ID>1919 </input>
<input>
<ID>IN_1</ID>1920 </input>
<input>
<ID>IN_2</ID>1921 </input>
<input>
<ID>IN_3</ID>1922 </input>
<input>
<ID>IN_B_0</ID>1941 </input>
<input>
<ID>IN_B_1</ID>1942 </input>
<input>
<ID>IN_B_2</ID>1939 </input>
<input>
<ID>IN_B_3</ID>1918 </input>
<output>
<ID>OUT_0</ID>1927 </output>
<output>
<ID>OUT_1</ID>1928 </output>
<output>
<ID>OUT_2</ID>1929 </output>
<output>
<ID>OUT_3</ID>1930 </output>
<output>
<ID>carry_out</ID>1913 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1329</ID>
<type>AE_FULLADDER_4BIT</type>
<position>668.5,1396</position>
<input>
<ID>IN_0</ID>1923 </input>
<input>
<ID>IN_1</ID>1924 </input>
<input>
<ID>IN_2</ID>1925 </input>
<input>
<ID>IN_3</ID>1926 </input>
<input>
<ID>IN_B_0</ID>1935 </input>
<input>
<ID>IN_B_1</ID>1936 </input>
<input>
<ID>IN_B_2</ID>1937 </input>
<input>
<ID>IN_B_3</ID>1938 </input>
<output>
<ID>OUT_0</ID>1931 </output>
<output>
<ID>OUT_1</ID>1932 </output>
<output>
<ID>OUT_2</ID>1933 </output>
<output>
<ID>OUT_3</ID>1934 </output>
<input>
<ID>carry_in</ID>1913 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1331</ID>
<type>DE_TO</type>
<position>709,1347</position>
<input>
<ID>IN_0</ID>1622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-3</lparam></gate>
<gate>
<ID>1332</ID>
<type>DE_TO</type>
<position>709,1337</position>
<input>
<ID>IN_0</ID>1664 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-4</lparam></gate>
<gate>
<ID>1333</ID>
<type>DE_TO</type>
<position>709,1335</position>
<input>
<ID>IN_0</ID>1783 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-5</lparam></gate>
<gate>
<ID>1334</ID>
<type>DA_FROM</type>
<position>662,1412.5</position>
<input>
<ID>IN_0</ID>1918 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1335</ID>
<type>DA_FROM</type>
<position>662,1388.5</position>
<input>
<ID>IN_0</ID>1926 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC7</lparam></gate>
<gate>
<ID>1336</ID>
<type>DA_FROM</type>
<position>662,1390.5</position>
<input>
<ID>IN_0</ID>1925 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC6</lparam></gate>
<gate>
<ID>1337</ID>
<type>DA_FROM</type>
<position>662,1392.5</position>
<input>
<ID>IN_0</ID>1924 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC5</lparam></gate>
<gate>
<ID>1338</ID>
<type>DA_FROM</type>
<position>662,1394.5</position>
<input>
<ID>IN_0</ID>1923 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC4</lparam></gate>
<gate>
<ID>1339</ID>
<type>DA_FROM</type>
<position>662,1406.5</position>
<input>
<ID>IN_0</ID>1921 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC2</lparam></gate>
<gate>
<ID>1340</ID>
<type>DA_FROM</type>
<position>662,1404.5</position>
<input>
<ID>IN_0</ID>1922 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC3</lparam></gate>
<gate>
<ID>1341</ID>
<type>DA_FROM</type>
<position>662,1408.5</position>
<input>
<ID>IN_0</ID>1920 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC1</lparam></gate>
<gate>
<ID>1342</ID>
<type>DA_FROM</type>
<position>662,1410.5</position>
<input>
<ID>IN_0</ID>1919 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC0</lparam></gate>
<gate>
<ID>1343</ID>
<type>DE_TO</type>
<position>675,1415</position>
<input>
<ID>IN_0</ID>1927 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-0</lparam></gate>
<gate>
<ID>1344</ID>
<type>DE_TO</type>
<position>675,1413</position>
<input>
<ID>IN_0</ID>1928 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-1</lparam></gate>
<gate>
<ID>1345</ID>
<type>DE_TO</type>
<position>675,1411</position>
<input>
<ID>IN_0</ID>1929 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-2</lparam></gate>
<gate>
<ID>1346</ID>
<type>DE_TO</type>
<position>675,1409</position>
<input>
<ID>IN_0</ID>1930 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-3</lparam></gate>
<gate>
<ID>1347</ID>
<type>DE_TO</type>
<position>675,1399</position>
<input>
<ID>IN_0</ID>1931 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-4</lparam></gate>
<gate>
<ID>1348</ID>
<type>DE_TO</type>
<position>675,1397</position>
<input>
<ID>IN_0</ID>1932 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-5</lparam></gate>
<gate>
<ID>1349</ID>
<type>DE_TO</type>
<position>675,1395</position>
<input>
<ID>IN_0</ID>1933 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-6</lparam></gate>
<gate>
<ID>1350</ID>
<type>DE_TO</type>
<position>675,1393</position>
<input>
<ID>IN_0</ID>1934 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-7</lparam></gate>
<gate>
<ID>1351</ID>
<type>DA_FROM</type>
<position>662,1402.5</position>
<input>
<ID>IN_0</ID>1935 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1352</ID>
<type>DA_FROM</type>
<position>662,1400.5</position>
<input>
<ID>IN_0</ID>1936 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1353</ID>
<type>DA_FROM</type>
<position>662,1398.5</position>
<input>
<ID>IN_0</ID>1937 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1354</ID>
<type>DA_FROM</type>
<position>662,1396.5</position>
<input>
<ID>IN_0</ID>1938 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1355</ID>
<type>DA_FROM</type>
<position>662,1414.5</position>
<input>
<ID>IN_0</ID>1939 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1356</ID>
<type>DE_TO</type>
<position>640.5,1390.5</position>
<input>
<ID>IN_0</ID>1940 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID off3sign</lparam></gate>
<gate>
<ID>1357</ID>
<type>DE_TO</type>
<position>709,1333</position>
<input>
<ID>IN_0</ID>1837 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-6</lparam></gate>
<gate>
<ID>1358</ID>
<type>BA_DECODER_2x4</type>
<position>628,1402</position>
<input>
<ID>ENABLE</ID>1949 </input>
<input>
<ID>IN_0</ID>1948 </input>
<output>
<ID>OUT_0</ID>1943 </output>
<output>
<ID>OUT_1</ID>1944 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1359</ID>
<type>DE_TO</type>
<position>709,1331</position>
<input>
<ID>IN_0</ID>1997 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-7</lparam></gate>
<gate>
<ID>1361</ID>
<type>EE_VDD</type>
<position>697,1356.5</position>
<output>
<ID>OUT_0</ID>1998 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1362</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>491.5,1383</position>
<input>
<ID>ENABLE_0</ID>2077 </input>
<input>
<ID>IN_0</ID>2046 </input>
<input>
<ID>IN_1</ID>2045 </input>
<input>
<ID>IN_2</ID>2044 </input>
<input>
<ID>IN_3</ID>2014 </input>
<input>
<ID>IN_4</ID>2008 </input>
<input>
<ID>IN_5</ID>2007 </input>
<input>
<ID>IN_6</ID>2000 </input>
<input>
<ID>IN_7</ID>1999 </input>
<output>
<ID>OUT_0</ID>2055 </output>
<output>
<ID>OUT_1</ID>2057 </output>
<output>
<ID>OUT_2</ID>2053 </output>
<output>
<ID>OUT_3</ID>2058 </output>
<output>
<ID>OUT_4</ID>2054 </output>
<output>
<ID>OUT_5</ID>2056 </output>
<output>
<ID>OUT_6</ID>2059 </output>
<output>
<ID>OUT_7</ID>2060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1363</ID>
<type>DA_FROM</type>
<position>479.5,1389.5</position>
<input>
<ID>IN_0</ID>1999 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-7</lparam></gate>
<gate>
<ID>1364</ID>
<type>DE_TO</type>
<position>661,1333</position>
<input>
<ID>IN_0</ID>1947 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BRop</lparam></gate>
<gate>
<ID>1365</ID>
<type>DA_FROM</type>
<position>479.5,1387.5</position>
<input>
<ID>IN_0</ID>2000 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-6</lparam></gate>
<gate>
<ID>1366</ID>
<type>DA_FROM</type>
<position>623,1400.5</position>
<input>
<ID>IN_0</ID>1948 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BR</lparam></gate>
<gate>
<ID>1367</ID>
<type>DA_FROM</type>
<position>479.5,1385.5</position>
<input>
<ID>IN_0</ID>2007 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-5</lparam></gate>
<gate>
<ID>1368</ID>
<type>AE_OR2</type>
<position>622,1403.5</position>
<input>
<ID>IN_0</ID>1952 </input>
<input>
<ID>IN_1</ID>1950 </input>
<output>
<ID>OUT</ID>1949 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1369</ID>
<type>DA_FROM</type>
<position>617,1402.5</position>
<input>
<ID>IN_0</ID>1950 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID BR</lparam></gate>
<gate>
<ID>1370</ID>
<type>DA_FROM</type>
<position>479.5,1383.5</position>
<input>
<ID>IN_0</ID>2008 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-4</lparam></gate>
<gate>
<ID>1371</ID>
<type>DE_TO</type>
<position>655,1353</position>
<input>
<ID>IN_0</ID>1951 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD/ST</lparam></gate>
<gate>
<ID>1372</ID>
<type>DA_FROM</type>
<position>479.5,1381.5</position>
<input>
<ID>IN_0</ID>2014 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-3</lparam></gate>
<gate>
<ID>1373</ID>
<type>DA_FROM</type>
<position>617,1404.5</position>
<input>
<ID>IN_0</ID>1952 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD/ST</lparam></gate>
<gate>
<ID>1374</ID>
<type>DA_FROM</type>
<position>479.5,1379.5</position>
<input>
<ID>IN_0</ID>2044 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-2</lparam></gate>
<gate>
<ID>1375</ID>
<type>DA_FROM</type>
<position>479.5,1377.5</position>
<input>
<ID>IN_0</ID>2045 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-1</lparam></gate>
<gate>
<ID>1376</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>491.5,1366</position>
<input>
<ID>ENABLE_0</ID>1962 </input>
<input>
<ID>IN_0</ID>1961 </input>
<input>
<ID>IN_1</ID>1960 </input>
<input>
<ID>IN_2</ID>1959 </input>
<input>
<ID>IN_3</ID>1958 </input>
<input>
<ID>IN_4</ID>1957 </input>
<input>
<ID>IN_5</ID>1956 </input>
<input>
<ID>IN_6</ID>1955 </input>
<input>
<ID>IN_7</ID>1954 </input>
<output>
<ID>OUT_0</ID>2055 </output>
<output>
<ID>OUT_1</ID>2057 </output>
<output>
<ID>OUT_2</ID>2053 </output>
<output>
<ID>OUT_3</ID>2058 </output>
<output>
<ID>OUT_4</ID>2054 </output>
<output>
<ID>OUT_5</ID>2056 </output>
<output>
<ID>OUT_6</ID>2059 </output>
<output>
<ID>OUT_7</ID>2060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1377</ID>
<type>DA_FROM</type>
<position>479.5,1373.5</position>
<input>
<ID>IN_0</ID>1954 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-7</lparam></gate>
<gate>
<ID>1378</ID>
<type>DA_FROM</type>
<position>479.5,1371.5</position>
<input>
<ID>IN_0</ID>1955 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-6</lparam></gate>
<gate>
<ID>1379</ID>
<type>DA_FROM</type>
<position>479.5,1369.5</position>
<input>
<ID>IN_0</ID>1956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-5</lparam></gate>
<gate>
<ID>1380</ID>
<type>DA_FROM</type>
<position>479.5,1367.5</position>
<input>
<ID>IN_0</ID>1957 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-4</lparam></gate>
<gate>
<ID>1381</ID>
<type>DA_FROM</type>
<position>479.5,1365.5</position>
<input>
<ID>IN_0</ID>1958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-3</lparam></gate>
<gate>
<ID>1382</ID>
<type>DA_FROM</type>
<position>479.5,1363.5</position>
<input>
<ID>IN_0</ID>1959 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-2</lparam></gate>
<gate>
<ID>1383</ID>
<type>DA_FROM</type>
<position>479.5,1361.5</position>
<input>
<ID>IN_0</ID>1960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-1</lparam></gate>
<gate>
<ID>1384</ID>
<type>DA_FROM</type>
<position>479.5,1359.5</position>
<input>
<ID>IN_0</ID>1961 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pcoff3-0</lparam></gate>
<gate>
<ID>1385</ID>
<type>DA_FROM</type>
<position>491.5,1373</position>
<input>
<ID>IN_0</ID>1962 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID BR</lparam></gate>
<gate>
<ID>1386</ID>
<type>DA_FROM</type>
<position>430,1384.5</position>
<input>
<ID>IN_0</ID>1963 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID LD/ST</lparam></gate>
<gate>
<ID>1387</ID>
<type>DA_FROM</type>
<position>479.5,1375.5</position>
<input>
<ID>IN_0</ID>2046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID pc+1-0</lparam></gate>
<gate>
<ID>1393</ID>
<type>AA_LABEL</type>
<position>667,1423</position>
<gparam>LABEL_TEXT PC + off3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1405</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>618,1337.5</position>
<input>
<ID>ENABLE_0</ID>2086 </input>
<input>
<ID>IN_0</ID>1642 </input>
<input>
<ID>IN_1</ID>1641 </input>
<input>
<ID>IN_2</ID>1640 </input>
<input>
<ID>IN_3</ID>1639 </input>
<input>
<ID>IN_4</ID>1638 </input>
<input>
<ID>IN_5</ID>1637 </input>
<input>
<ID>IN_6</ID>1636 </input>
<input>
<ID>IN_7</ID>1635 </input>
<output>
<ID>OUT_0</ID>1976 </output>
<output>
<ID>OUT_1</ID>1977 </output>
<output>
<ID>OUT_2</ID>1978 </output>
<output>
<ID>OUT_3</ID>1979 </output>
<output>
<ID>OUT_4</ID>1980 </output>
<output>
<ID>OUT_5</ID>1981 </output>
<output>
<ID>OUT_6</ID>1982 </output>
<output>
<ID>OUT_7</ID>1983 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1406</ID>
<type>AE_SMALL_INVERTER</type>
<position>491.5,1390</position>
<input>
<ID>IN_0</ID>2052 </input>
<output>
<ID>OUT_0</ID>2077 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1409</ID>
<type>DE_TO</type>
<position>631.5,1327</position>
<input>
<ID>IN_0</ID>1976 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr0</lparam></gate>
<gate>
<ID>1410</ID>
<type>DE_TO</type>
<position>631.5,1329</position>
<input>
<ID>IN_0</ID>1977 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr1</lparam></gate>
<gate>
<ID>1411</ID>
<type>DA_FROM</type>
<position>491.5,1394</position>
<input>
<ID>IN_0</ID>2052 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID BR</lparam></gate>
<gate>
<ID>1412</ID>
<type>EE_VDD</type>
<position>532,1319.5</position>
<output>
<ID>OUT_0</ID>1519 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1413</ID>
<type>DE_TO</type>
<position>631.5,1331</position>
<input>
<ID>IN_0</ID>1978 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr2</lparam></gate>
<gate>
<ID>1414</ID>
<type>DE_TO</type>
<position>631.5,1333</position>
<input>
<ID>IN_0</ID>1979 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr3</lparam></gate>
<gate>
<ID>1415</ID>
<type>DE_TO</type>
<position>631.5,1335</position>
<input>
<ID>IN_0</ID>1980 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr4</lparam></gate>
<gate>
<ID>1416</ID>
<type>DE_TO</type>
<position>631.5,1337</position>
<input>
<ID>IN_0</ID>1981 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr5</lparam></gate>
<gate>
<ID>1417</ID>
<type>DE_TO</type>
<position>631.5,1339</position>
<input>
<ID>IN_0</ID>1982 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr6</lparam></gate>
<gate>
<ID>1418</ID>
<type>DE_TO</type>
<position>631.5,1341</position>
<input>
<ID>IN_0</ID>1983 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr7</lparam></gate>
<gate>
<ID>1420</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>509,1326.5</position>
<input>
<ID>ENABLE_0</ID>1846 </input>
<input>
<ID>IN_0</ID>1760 </input>
<input>
<ID>IN_1</ID>1759 </input>
<input>
<ID>IN_2</ID>1758 </input>
<input>
<ID>IN_3</ID>1757 </input>
<input>
<ID>IN_4</ID>1756 </input>
<input>
<ID>IN_5</ID>1755 </input>
<input>
<ID>IN_6</ID>1754 </input>
<input>
<ID>IN_7</ID>1753 </input>
<output>
<ID>OUT_0</ID>1847 </output>
<output>
<ID>OUT_1</ID>1915 </output>
<output>
<ID>OUT_2</ID>1916 </output>
<output>
<ID>OUT_3</ID>1914 </output>
<output>
<ID>OUT_4</ID>1875 </output>
<output>
<ID>OUT_5</ID>1894 </output>
<output>
<ID>OUT_6</ID>1912 </output>
<output>
<ID>OUT_7</ID>1857 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1422</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>617.5,1348.5</position>
<input>
<ID>ENABLE_0</ID>2087 </input>
<input>
<ID>IN_0</ID>1642 </input>
<input>
<ID>IN_1</ID>1641 </input>
<input>
<ID>IN_2</ID>1640 </input>
<input>
<ID>IN_3</ID>1639 </input>
<input>
<ID>IN_4</ID>1638 </input>
<input>
<ID>IN_5</ID>1637 </input>
<input>
<ID>IN_6</ID>1636 </input>
<input>
<ID>IN_7</ID>1635 </input>
<output>
<ID>OUT_0</ID>2064 </output>
<output>
<ID>OUT_1</ID>2068 </output>
<output>
<ID>OUT_2</ID>2067 </output>
<output>
<ID>OUT_3</ID>2065 </output>
<output>
<ID>OUT_4</ID>2063 </output>
<output>
<ID>OUT_5</ID>2066 </output>
<output>
<ID>OUT_6</ID>2069 </output>
<output>
<ID>OUT_7</ID>2062 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1423</ID>
<type>DA_FROM</type>
<position>392.5,1267</position>
<input>
<ID>IN_0</ID>1984 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr0</lparam></gate>
<gate>
<ID>1424</ID>
<type>DA_FROM</type>
<position>392.5,1269</position>
<input>
<ID>IN_0</ID>1991 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr1</lparam></gate>
<gate>
<ID>1425</ID>
<type>DA_FROM</type>
<position>392.5,1271</position>
<input>
<ID>IN_0</ID>1990 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr2</lparam></gate>
<gate>
<ID>1426</ID>
<type>DA_FROM</type>
<position>392.5,1273</position>
<input>
<ID>IN_0</ID>1989 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr3</lparam></gate>
<gate>
<ID>1427</ID>
<type>DA_FROM</type>
<position>392.5,1275</position>
<input>
<ID>IN_0</ID>1988 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr4</lparam></gate>
<gate>
<ID>1428</ID>
<type>DA_FROM</type>
<position>392.5,1277</position>
<input>
<ID>IN_0</ID>1987 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr5</lparam></gate>
<gate>
<ID>1429</ID>
<type>DA_FROM</type>
<position>392.5,1279</position>
<input>
<ID>IN_0</ID>1986 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr6</lparam></gate>
<gate>
<ID>1430</ID>
<type>DA_FROM</type>
<position>392.5,1281</position>
<input>
<ID>IN_0</ID>1985 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr7</lparam></gate>
<gate>
<ID>1435</ID>
<type>DA_FROM</type>
<position>505.5,1332.5</position>
<input>
<ID>IN_0</ID>1846 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>1438</ID>
<type>EE_VDD</type>
<position>607,1355</position>
<output>
<ID>OUT_0</ID>2072 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1439</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>591.5,1338.5</position>
<input>
<ID>ENABLE_0</ID>1917 </input>
<input>
<ID>IN_0</ID>1847 </input>
<input>
<ID>IN_1</ID>1915 </input>
<input>
<ID>IN_2</ID>1916 </input>
<input>
<ID>IN_3</ID>1914 </input>
<input>
<ID>IN_4</ID>1875 </input>
<input>
<ID>IN_5</ID>1894 </input>
<input>
<ID>IN_6</ID>1912 </input>
<input>
<ID>IN_7</ID>1857 </input>
<output>
<ID>OUT_0</ID>1654 </output>
<output>
<ID>OUT_1</ID>1655 </output>
<output>
<ID>OUT_2</ID>1656 </output>
<output>
<ID>OUT_3</ID>1657 </output>
<output>
<ID>OUT_4</ID>1658 </output>
<output>
<ID>OUT_5</ID>1653 </output>
<output>
<ID>OUT_6</ID>1660 </output>
<output>
<ID>OUT_7</ID>1659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1440</ID>
<type>DA_FROM</type>
<position>588.5,1343.5</position>
<input>
<ID>IN_0</ID>1917 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>1454</ID>
<type>DA_FROM</type>
<position>553,1354</position>
<input>
<ID>IN_0</ID>1995 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>1455</ID>
<type>DA_FROM</type>
<position>422.5,1312.5</position>
<input>
<ID>IN_0</ID>1996 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD</lparam></gate>
<gate>
<ID>1457</ID>
<type>DA_FROM</type>
<position>595,1393</position>
<input>
<ID>IN_0</ID>1645 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>1466</ID>
<type>DA_FROM</type>
<position>399.5,1332</position>
<input>
<ID>IN_0</ID>2001 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STR</lparam></gate>
<gate>
<ID>1467</ID>
<type>DA_FROM</type>
<position>407.5,1285</position>
<input>
<ID>IN_0</ID>2002 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD</lparam></gate>
<gate>
<ID>1469</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>413.5,1265</position>
<input>
<ID>ENABLE_0</ID>2003 </input>
<input>
<ID>IN_0</ID>2022 </input>
<input>
<ID>IN_1</ID>2021 </input>
<input>
<ID>IN_2</ID>2020 </input>
<input>
<ID>IN_3</ID>2019 </input>
<input>
<ID>IN_4</ID>2018 </input>
<input>
<ID>IN_5</ID>2017 </input>
<input>
<ID>IN_6</ID>2016 </input>
<input>
<ID>IN_7</ID>2015 </input>
<output>
<ID>OUT_0</ID>1782 </output>
<output>
<ID>OUT_1</ID>1781 </output>
<output>
<ID>OUT_2</ID>1780 </output>
<output>
<ID>OUT_3</ID>1779 </output>
<output>
<ID>OUT_4</ID>1778 </output>
<output>
<ID>OUT_5</ID>1777 </output>
<output>
<ID>OUT_6</ID>1776 </output>
<output>
<ID>OUT_7</ID>1775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1471</ID>
<type>EE_VDD</type>
<position>413.5,1271.5</position>
<output>
<ID>OUT_0</ID>2003 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1479</ID>
<type>EE_VDD</type>
<position>618,1343.5</position>
<output>
<ID>OUT_0</ID>2086 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1481</ID>
<type>EE_VDD</type>
<position>617.5,1354.5</position>
<output>
<ID>OUT_0</ID>2087 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1483</ID>
<type>AA_TOGGLE</type>
<position>622,1355.5</position>
<output>
<ID>OUT_0</ID>2088 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1485</ID>
<type>DA_FROM</type>
<position>404,1254.5</position>
<input>
<ID>IN_0</ID>2022 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU0</lparam></gate>
<gate>
<ID>1486</ID>
<type>DA_FROM</type>
<position>404,1256.5</position>
<input>
<ID>IN_0</ID>2021 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU1</lparam></gate>
<gate>
<ID>1487</ID>
<type>DA_FROM</type>
<position>404,1258.5</position>
<input>
<ID>IN_0</ID>2020 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU2</lparam></gate>
<gate>
<ID>1488</ID>
<type>DA_FROM</type>
<position>404,1260.5</position>
<input>
<ID>IN_0</ID>2019 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU3</lparam></gate>
<gate>
<ID>1489</ID>
<type>DA_FROM</type>
<position>404,1262.5</position>
<input>
<ID>IN_0</ID>2018 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU4</lparam></gate>
<gate>
<ID>1490</ID>
<type>DA_FROM</type>
<position>404,1264.5</position>
<input>
<ID>IN_0</ID>2017 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU5</lparam></gate>
<gate>
<ID>1491</ID>
<type>DA_FROM</type>
<position>404,1266.5</position>
<input>
<ID>IN_0</ID>2016 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU6</lparam></gate>
<gate>
<ID>1492</ID>
<type>DA_FROM</type>
<position>404,1268.5</position>
<input>
<ID>IN_0</ID>2015 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU7</lparam></gate>
<gate>
<ID>1493</ID>
<type>AE_SMALL_INVERTER</type>
<position>430,1369.5</position>
<input>
<ID>IN_0</ID>2076 </input>
<output>
<ID>OUT_0</ID>2090 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1494</ID>
<type>DA_FROM</type>
<position>568,1330</position>
<input>
<ID>IN_0</ID>1665 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>1496</ID>
<type>EE_VDD</type>
<position>573.5,1332.5</position>
<output>
<ID>OUT_0</ID>2023 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1498</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>404,1317</position>
<input>
<ID>ENABLE_0</ID>2024 </input>
<input>
<ID>IN_0</ID>2032 </input>
<input>
<ID>IN_1</ID>2031 </input>
<input>
<ID>IN_2</ID>2030 </input>
<input>
<ID>IN_3</ID>2029 </input>
<output>
<ID>OUT_0</ID>1763 </output>
<output>
<ID>OUT_1</ID>1764 </output>
<output>
<ID>OUT_2</ID>1773 </output>
<output>
<ID>OUT_3</ID>1774 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1500</ID>
<type>AE_OR2</type>
<position>408,1301</position>
<input>
<ID>IN_0</ID>2025 </input>
<input>
<ID>IN_1</ID>2026 </input>
<output>
<ID>OUT</ID>2024 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1501</ID>
<type>AA_LABEL</type>
<position>563,1429</position>
<gparam>LABEL_TEXT GWLC</gparam>
<gparam>TEXT_HEIGHT 20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1502</ID>
<type>DA_FROM</type>
<position>403,1302</position>
<input>
<ID>IN_0</ID>2025 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>1504</ID>
<type>DA_FROM</type>
<position>403,1300</position>
<input>
<ID>IN_0</ID>2026 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>1505</ID>
<type>AA_LABEL</type>
<position>654,1286.5</position>
<gparam>LABEL_TEXT Easy to read ADD output</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1506</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>427.5,1298</position>
<input>
<ID>ENABLE_0</ID>2024 </input>
<input>
<ID>IN_0</ID>2028 </input>
<input>
<ID>IN_1</ID>2027 </input>
<output>
<ID>OUT_0</ID>1601 </output>
<output>
<ID>OUT_1</ID>1600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1507</ID>
<type>DA_FROM</type>
<position>422,1298</position>
<input>
<ID>IN_0</ID>2027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr5</lparam></gate>
<gate>
<ID>1508</ID>
<type>DA_FROM</type>
<position>422,1296</position>
<input>
<ID>IN_0</ID>2028 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr4</lparam></gate>
<gate>
<ID>1509</ID>
<type>DA_FROM</type>
<position>397.5,1312.5</position>
<input>
<ID>IN_0</ID>2032 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr0</lparam></gate>
<gate>
<ID>1510</ID>
<type>DA_FROM</type>
<position>397.5,1314.5</position>
<input>
<ID>IN_0</ID>2031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr1</lparam></gate>
<gate>
<ID>1511</ID>
<type>DA_FROM</type>
<position>397.5,1316.5</position>
<input>
<ID>IN_0</ID>2030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr2</lparam></gate>
<gate>
<ID>1512</ID>
<type>DA_FROM</type>
<position>397.5,1318.5</position>
<input>
<ID>IN_0</ID>2029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mdr3</lparam></gate>
<gate>
<ID>1513</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>671.5,1279.5</position>
<input>
<ID>ENABLE_0</ID>2041 </input>
<input>
<ID>IN_0</ID>1717 </input>
<input>
<ID>IN_1</ID>1718 </input>
<input>
<ID>IN_2</ID>1719 </input>
<input>
<ID>IN_3</ID>1720 </input>
<input>
<ID>IN_4</ID>1721 </input>
<input>
<ID>IN_5</ID>1722 </input>
<input>
<ID>IN_6</ID>1723 </input>
<input>
<ID>IN_7</ID>1724 </input>
<output>
<ID>OUT_0</ID>2040 </output>
<output>
<ID>OUT_1</ID>2039 </output>
<output>
<ID>OUT_2</ID>2038 </output>
<output>
<ID>OUT_3</ID>2035 </output>
<output>
<ID>OUT_4</ID>2037 </output>
<output>
<ID>OUT_5</ID>2034 </output>
<output>
<ID>OUT_6</ID>2036 </output>
<output>
<ID>OUT_7</ID>2033 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1514</ID>
<type>DE_TO</type>
<position>695,1283</position>
<input>
<ID>IN_0</ID>2033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU7</lparam></gate>
<gate>
<ID>1515</ID>
<type>DE_TO</type>
<position>695,1281</position>
<input>
<ID>IN_0</ID>2034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU5</lparam></gate>
<gate>
<ID>1516</ID>
<type>DE_TO</type>
<position>695,1279</position>
<input>
<ID>IN_0</ID>2035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU3</lparam></gate>
<gate>
<ID>1517</ID>
<type>DE_TO</type>
<position>703,1282</position>
<input>
<ID>IN_0</ID>2036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU6</lparam></gate>
<gate>
<ID>1518</ID>
<type>DE_TO</type>
<position>703,1280</position>
<input>
<ID>IN_0</ID>2037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU4</lparam></gate>
<gate>
<ID>1519</ID>
<type>DE_TO</type>
<position>703,1278</position>
<input>
<ID>IN_0</ID>2038 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU2</lparam></gate>
<gate>
<ID>1520</ID>
<type>DE_TO</type>
<position>695,1277</position>
<input>
<ID>IN_0</ID>2039 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU1</lparam></gate>
<gate>
<ID>1521</ID>
<type>DE_TO</type>
<position>703,1276</position>
<input>
<ID>IN_0</ID>2040 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU0</lparam></gate>
<gate>
<ID>1523</ID>
<type>AA_LABEL</type>
<position>622,1358</position>
<gparam>LABEL_TEXT IR Load Control</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1525</ID>
<type>AE_OR2</type>
<position>671.5,1287.5</position>
<input>
<ID>IN_0</ID>2042 </input>
<input>
<ID>IN_1</ID>2043 </input>
<output>
<ID>OUT</ID>2041 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1526</ID>
<type>AA_LABEL</type>
<position>507.5,1384</position>
<gparam>LABEL_TEXT PC INPUT</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1527</ID>
<type>DA_FROM</type>
<position>672.5,1292.5</position>
<input>
<ID>IN_0</ID>2042 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>1528</ID>
<type>DA_FROM</type>
<position>670.5,1292.5</position>
<input>
<ID>IN_0</ID>2043 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>1530</ID>
<type>AA_LABEL</type>
<position>415,1329.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1532</ID>
<type>AE_OR3</type>
<position>410,1340.5</position>
<input>
<ID>IN_0</ID>2070 </input>
<input>
<ID>IN_1</ID>2071 </input>
<input>
<ID>IN_2</ID>2073 </input>
<output>
<ID>OUT</ID>2074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1534</ID>
<type>DA_FROM</type>
<position>405,1342.5</position>
<input>
<ID>IN_0</ID>2070 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LD</lparam></gate>
<gate>
<ID>1536</ID>
<type>DA_FROM</type>
<position>405,1340.5</position>
<input>
<ID>IN_0</ID>2071 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<wire>
<ID>1553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697.5,1343.5,697.5,1345</points>
<intersection>1343.5 4</intersection>
<intersection>1345 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>697.5,1345,698.5,1345</points>
<connection>
<GID>1177</GID>
<name>IN_3</name></connection>
<intersection>697.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>697.5,1343.5,698,1343.5</points>
<connection>
<GID>1297</GID>
<name>IN_0</name></connection>
<intersection>697.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1554</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>663.5,1356,663.5,1357.5</points>
<connection>
<GID>1055</GID>
<name>OUT_0</name></connection>
<intersection>1356 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>663.5,1356,665,1356</points>
<connection>
<GID>965</GID>
<name>IN_1</name></connection>
<intersection>663.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1555</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>653,1337.5,653,1341</points>
<connection>
<GID>1052</GID>
<name>IN_1</name></connection>
<connection>
<GID>1071</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457,1287.5,485,1287.5</points>
<connection>
<GID>1145</GID>
<name>IN_3</name></connection>
<connection>
<GID>1166</GID>
<name>IN_3</name></connection>
<intersection>457 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>457,1286.5,457,1287.5</points>
<intersection>1286.5 8</intersection>
<intersection>1287.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>454,1286.5,457,1286.5</points>
<connection>
<GID>1103</GID>
<name>OUT_2</name></connection>
<intersection>457 7</intersection></hsegment></shape></wire>
<wire>
<ID>1557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524,1379.5,524,1391.5</points>
<intersection>1379.5 2</intersection>
<intersection>1383.5 4</intersection>
<intersection>1391.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>523,1379.5,524,1379.5</points>
<connection>
<GID>1063</GID>
<name>OUT_0</name></connection>
<intersection>524 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1391.5,524,1391.5</points>
<connection>
<GID>1061</GID>
<name>OUT_0</name></connection>
<intersection>524 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>524,1383.5,532,1383.5</points>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection>
<intersection>524 0</intersection></hsegment></shape></wire>
<wire>
<ID>1558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>524.5,1380.5,524.5,1392.5</points>
<intersection>1380.5 2</intersection>
<intersection>1384.5 1</intersection>
<intersection>1392.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>524.5,1384.5,532,1384.5</points>
<connection>
<GID>1065</GID>
<name>IN_1</name></connection>
<intersection>524.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>523,1380.5,524.5,1380.5</points>
<connection>
<GID>1063</GID>
<name>OUT_1</name></connection>
<intersection>524.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1392.5,524.5,1392.5</points>
<connection>
<GID>1061</GID>
<name>OUT_1</name></connection>
<intersection>524.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525,1381.5,525,1393.5</points>
<intersection>1381.5 2</intersection>
<intersection>1385.5 1</intersection>
<intersection>1393.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1385.5,532,1385.5</points>
<connection>
<GID>1065</GID>
<name>IN_2</name></connection>
<intersection>525 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>523,1381.5,525,1381.5</points>
<connection>
<GID>1063</GID>
<name>OUT_2</name></connection>
<intersection>525 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1393.5,525,1393.5</points>
<connection>
<GID>1061</GID>
<name>OUT_2</name></connection>
<intersection>525 0</intersection></hsegment></shape></wire>
<wire>
<ID>1560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525.5,1382.5,525.5,1394.5</points>
<intersection>1382.5 1</intersection>
<intersection>1386.5 2</intersection>
<intersection>1394.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>523,1382.5,525.5,1382.5</points>
<connection>
<GID>1063</GID>
<name>OUT_3</name></connection>
<intersection>525.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525.5,1386.5,532,1386.5</points>
<connection>
<GID>1065</GID>
<name>IN_3</name></connection>
<intersection>525.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1394.5,525.5,1394.5</points>
<connection>
<GID>1061</GID>
<name>OUT_3</name></connection>
<intersection>525.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>526,1383.5,526,1395.5</points>
<intersection>1383.5 1</intersection>
<intersection>1387.5 5</intersection>
<intersection>1395.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>523,1383.5,526,1383.5</points>
<connection>
<GID>1063</GID>
<name>OUT_4</name></connection>
<intersection>526 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1395.5,526,1395.5</points>
<connection>
<GID>1061</GID>
<name>OUT_4</name></connection>
<intersection>526 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>526,1387.5,532,1387.5</points>
<connection>
<GID>1065</GID>
<name>IN_4</name></connection>
<intersection>526 0</intersection></hsegment></shape></wire>
<wire>
<ID>1562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>526.5,1384.5,526.5,1396.5</points>
<intersection>1384.5 1</intersection>
<intersection>1388.5 2</intersection>
<intersection>1396.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>523,1384.5,526.5,1384.5</points>
<connection>
<GID>1063</GID>
<name>OUT_5</name></connection>
<intersection>526.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>526.5,1388.5,532,1388.5</points>
<connection>
<GID>1065</GID>
<name>IN_5</name></connection>
<intersection>526.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1396.5,526.5,1396.5</points>
<connection>
<GID>1061</GID>
<name>OUT_5</name></connection>
<intersection>526.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527,1385.5,527,1397.5</points>
<intersection>1385.5 1</intersection>
<intersection>1389.5 2</intersection>
<intersection>1397.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>523,1385.5,527,1385.5</points>
<connection>
<GID>1063</GID>
<name>OUT_6</name></connection>
<intersection>527 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527,1389.5,532,1389.5</points>
<connection>
<GID>1065</GID>
<name>IN_6</name></connection>
<intersection>527 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1397.5,527,1397.5</points>
<connection>
<GID>1061</GID>
<name>OUT_6</name></connection>
<intersection>527 0</intersection></hsegment></shape></wire>
<wire>
<ID>1564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>527.5,1386.5,527.5,1398.5</points>
<intersection>1386.5 1</intersection>
<intersection>1390.5 2</intersection>
<intersection>1398.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>523,1386.5,527.5,1386.5</points>
<connection>
<GID>1063</GID>
<name>OUT_7</name></connection>
<intersection>527.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>527.5,1390.5,532,1390.5</points>
<connection>
<GID>1065</GID>
<name>IN_7</name></connection>
<intersection>527.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>523,1398.5,527.5,1398.5</points>
<connection>
<GID>1061</GID>
<name>OUT_7</name></connection>
<intersection>527.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513,1405.5,513,1407</points>
<connection>
<GID>1067</GID>
<name>ENABLE</name></connection>
<connection>
<GID>1069</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1566</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>512.5,1402.5,513,1402.5</points>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection>
<connection>
<GID>1072</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521,1388,521,1403</points>
<connection>
<GID>1063</GID>
<name>ENABLE_0</name></connection>
<intersection>1403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520,1403,521,1403</points>
<intersection>520 2</intersection>
<intersection>521 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>520,1402.5,520,1403</points>
<intersection>1402.5 3</intersection>
<intersection>1403 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>519,1402.5,520,1402.5</points>
<connection>
<GID>1067</GID>
<name>OUT_0</name></connection>
<intersection>520 2</intersection></hsegment></shape></wire>
<wire>
<ID>1568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521,1400,521,1403</points>
<connection>
<GID>1061</GID>
<name>ENABLE_0</name></connection>
<intersection>1403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520,1403,521,1403</points>
<intersection>520 2</intersection>
<intersection>521 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>520,1403,520,1403.5</points>
<intersection>1403 1</intersection>
<intersection>1403.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>519,1403.5,520,1403.5</points>
<connection>
<GID>1067</GID>
<name>OUT_1</name></connection>
<intersection>520 2</intersection></hsegment></shape></wire>
<wire>
<ID>1569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503,1391.5,503,1394</points>
<connection>
<GID>1074</GID>
<name>OUT_0</name></connection>
<intersection>1391.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503,1391.5,519,1391.5</points>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection>
<intersection>503 0</intersection></hsegment></shape></wire>
<wire>
<ID>1570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>503.5,1392.5,503.5,1396</points>
<intersection>1392.5 1</intersection>
<intersection>1396 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>503.5,1392.5,519,1392.5</points>
<connection>
<GID>1061</GID>
<name>IN_1</name></connection>
<intersection>503.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>503,1396,503.5,1396</points>
<connection>
<GID>1074</GID>
<name>OUT_1</name></connection>
<intersection>503.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504,1393.5,504,1398</points>
<intersection>1393.5 2</intersection>
<intersection>1398 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>504,1393.5,519,1393.5</points>
<connection>
<GID>1061</GID>
<name>IN_2</name></connection>
<intersection>504 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>503,1398,504,1398</points>
<connection>
<GID>1074</GID>
<name>OUT_2</name></connection>
<intersection>504 0</intersection></hsegment></shape></wire>
<wire>
<ID>1572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>504.5,1394.5,504.5,1400</points>
<intersection>1394.5 1</intersection>
<intersection>1400 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>504.5,1394.5,519,1394.5</points>
<connection>
<GID>1061</GID>
<name>IN_3</name></connection>
<intersection>504.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,1400,504.5,1400</points>
<connection>
<GID>1074</GID>
<name>OUT_3</name></connection>
<intersection>504.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505,1395.5,505,1406.5</points>
<intersection>1395.5 1</intersection>
<intersection>1406.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505,1395.5,519,1395.5</points>
<connection>
<GID>1061</GID>
<name>IN_4</name></connection>
<intersection>505 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,1406.5,505,1406.5</points>
<connection>
<GID>1073</GID>
<name>OUT_0</name></connection>
<intersection>505 0</intersection></hsegment></shape></wire>
<wire>
<ID>1574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,1396.5,505.5,1408.5</points>
<intersection>1396.5 1</intersection>
<intersection>1408.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505.5,1396.5,519,1396.5</points>
<connection>
<GID>1061</GID>
<name>IN_5</name></connection>
<intersection>505.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,1408.5,505.5,1408.5</points>
<connection>
<GID>1073</GID>
<name>OUT_1</name></connection>
<intersection>505.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506,1397.5,506,1410.5</points>
<intersection>1397.5 1</intersection>
<intersection>1410.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>506,1397.5,519,1397.5</points>
<connection>
<GID>1061</GID>
<name>IN_6</name></connection>
<intersection>506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,1410.5,506,1410.5</points>
<connection>
<GID>1073</GID>
<name>OUT_2</name></connection>
<intersection>506 0</intersection></hsegment></shape></wire>
<wire>
<ID>1576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>506.5,1398.5,506.5,1412.5</points>
<intersection>1398.5 1</intersection>
<intersection>1412.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>506.5,1398.5,519,1398.5</points>
<connection>
<GID>1061</GID>
<name>IN_7</name></connection>
<intersection>506.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>503,1412.5,506.5,1412.5</points>
<connection>
<GID>1073</GID>
<name>OUT_3</name></connection>
<intersection>506.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1389.5,545,1389.5</points>
<connection>
<GID>1102</GID>
<name>IN_6</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1388.5,545,1388.5</points>
<connection>
<GID>1102</GID>
<name>IN_5</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1383.5,545,1383.5</points>
<connection>
<GID>1102</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1390.5,545,1390.5</points>
<connection>
<GID>1102</GID>
<name>IN_7</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1581</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1386.5,545,1386.5</points>
<connection>
<GID>1102</GID>
<name>IN_3</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1384.5,545,1384.5</points>
<connection>
<GID>1102</GID>
<name>IN_1</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1385.5,545,1385.5</points>
<connection>
<GID>1102</GID>
<name>IN_2</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1387.5,545,1387.5</points>
<connection>
<GID>1102</GID>
<name>IN_4</name></connection>
<connection>
<GID>1065</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1586</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>468.5,1292.5,468.5,1327</points>
<intersection>1292.5 6</intersection>
<intersection>1327 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1327,468.5,1327</points>
<connection>
<GID>1138</GID>
<name>OUT_3</name></connection>
<intersection>468.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>468.5,1292.5,485,1292.5</points>
<connection>
<GID>1165</GID>
<name>IN_0</name></connection>
<connection>
<GID>1144</GID>
<name>IN_0</name></connection>
<intersection>468.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639,1334,639,1354</points>
<intersection>1334 6</intersection>
<intersection>1339.5 2</intersection>
<intersection>1345 11</intersection>
<intersection>1352 1</intersection>
<intersection>1354 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>629.5,1352,639,1352</points>
<connection>
<GID>1108</GID>
<name>OUT_7</name></connection>
<intersection>639 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639,1339.5,653,1339.5</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<intersection>639 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>639,1334,653,1334</points>
<connection>
<GID>1053</GID>
<name>IN_0</name></connection>
<intersection>639 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>639,1354,641.5,1354</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<intersection>639 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>639,1345,649,1345</points>
<connection>
<GID>1077</GID>
<name>IN_0</name></connection>
<intersection>639 0</intersection></hsegment></shape></wire>
<wire>
<ID>1595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>711.5,1290.5,711.5,1293</points>
<connection>
<GID>1075</GID>
<name>IN_0</name></connection>
<intersection>1290.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>711,1290.5,711.5,1290.5</points>
<connection>
<GID>1060</GID>
<name>OUT</name></connection>
<intersection>711.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,1333,448,1341</points>
<intersection>1333 2</intersection>
<intersection>1341 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,1341,448,1341</points>
<connection>
<GID>1181</GID>
<name>OUT_0</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,1333,449,1333</points>
<connection>
<GID>1138</GID>
<name>load</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>1597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,1320,448,1342</points>
<intersection>1320 2</intersection>
<intersection>1342 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,1342,448,1342</points>
<connection>
<GID>1181</GID>
<name>OUT_1</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,1320,449,1320</points>
<connection>
<GID>1136</GID>
<name>load</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>1598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,1306.5,448,1343</points>
<intersection>1306.5 2</intersection>
<intersection>1343 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,1343,448,1343</points>
<connection>
<GID>1181</GID>
<name>OUT_2</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,1306.5,449,1306.5</points>
<connection>
<GID>1105</GID>
<name>load</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>1599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,1293.5,448,1344</points>
<intersection>1293.5 2</intersection>
<intersection>1344 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,1344,448,1344</points>
<connection>
<GID>1181</GID>
<name>OUT_3</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>448,1293.5,449,1293.5</points>
<connection>
<GID>1103</GID>
<name>load</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>1600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,1297.5,431.5,1342</points>
<intersection>1297.5 6</intersection>
<intersection>1309 10</intersection>
<intersection>1342 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,1342,432,1342</points>
<connection>
<GID>1181</GID>
<name>IN_1</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>429.5,1297.5,431.5,1297.5</points>
<connection>
<GID>1506</GID>
<name>OUT_1</name></connection>
<intersection>431.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>429,1309,431.5,1309</points>
<connection>
<GID>1298</GID>
<name>OUT_1</name></connection>
<intersection>431.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,1296.5,432,1341</points>
<connection>
<GID>1181</GID>
<name>IN_0</name></connection>
<intersection>1296.5 12</intersection>
<intersection>1308 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>429,1308,432,1308</points>
<connection>
<GID>1298</GID>
<name>OUT_0</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>429.5,1296.5,432,1296.5</points>
<connection>
<GID>1506</GID>
<name>OUT_0</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>1602</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>698,1332,698,1333.5</points>
<connection>
<GID>1288</GID>
<name>IN_0</name></connection>
<intersection>1332 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>698,1332,698.5,1332</points>
<connection>
<GID>1179</GID>
<name>IN_0</name></connection>
<intersection>698 2</intersection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>671,1357,671.5,1357</points>
<connection>
<GID>965</GID>
<name>OUT</name></connection>
<connection>
<GID>967</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1603</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>698,1331.5,698.5,1331.5</points>
<connection>
<GID>1285</GID>
<name>IN_0</name></connection>
<intersection>698.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>698.5,1331,698.5,1331.5</points>
<connection>
<GID>1179</GID>
<name>IN_1</name></connection>
<intersection>1331.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>1604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522.5,1375,540.5,1375</points>
<connection>
<GID>1129</GID>
<name>IN_0</name></connection>
<connection>
<GID>1132</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>653,1345,653,1345</points>
<connection>
<GID>1077</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1296</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>639.5,1332,639.5,1352</points>
<intersection>1332 2</intersection>
<intersection>1341 3</intersection>
<intersection>1343 4</intersection>
<intersection>1351 1</intersection>
<intersection>1352 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>629.5,1351,639.5,1351</points>
<connection>
<GID>1108</GID>
<name>OUT_6</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>639.5,1332,653,1332</points>
<connection>
<GID>1053</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>639.5,1341,649,1341</points>
<connection>
<GID>1071</GID>
<name>IN_0</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>639.5,1343,653,1343</points>
<connection>
<GID>1296</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>639.5,1352,641.5,1352</points>
<connection>
<GID>1054</GID>
<name>IN_1</name></connection>
<intersection>639.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1607</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>717.5,1293,722.5,1293</points>
<connection>
<GID>1084</GID>
<name>IN_0</name></connection>
<connection>
<GID>1075</GID>
<name>OUT_0</name></connection>
<intersection>721 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>721,1293,721,1312.5</points>
<intersection>1293 1</intersection>
<intersection>1312.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>721,1312.5,734,1312.5</points>
<connection>
<GID>1028</GID>
<name>IN_1</name></connection>
<intersection>721 8</intersection></hsegment></shape></wire>
<wire>
<ID>1608</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>698.5,1329.5,698.5,1330</points>
<connection>
<GID>1179</GID>
<name>IN_2</name></connection>
<intersection>1329.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>698,1329.5,698.5,1329.5</points>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection>
<intersection>698.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1609</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>698.5,1327.5,698.5,1329</points>
<connection>
<GID>1179</GID>
<name>IN_3</name></connection>
<intersection>1327.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>698,1327.5,698.5,1327.5</points>
<connection>
<GID>1246</GID>
<name>IN_0</name></connection>
<intersection>698.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1610</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>717.5,1294,722.5,1294</points>
<connection>
<GID>1084</GID>
<name>IN_1</name></connection>
<connection>
<GID>1075</GID>
<name>OUT_1</name></connection>
<intersection>720.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>720.5,1294,720.5,1316.5</points>
<intersection>1294 1</intersection>
<intersection>1316.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>720.5,1316.5,734,1316.5</points>
<connection>
<GID>1026</GID>
<name>IN_1</name></connection>
<intersection>720.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1611</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>717.5,1295,722.5,1295</points>
<connection>
<GID>1084</GID>
<name>IN_2</name></connection>
<connection>
<GID>1075</GID>
<name>OUT_2</name></connection>
<intersection>720 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>720,1295,720,1320.5</points>
<intersection>1295 1</intersection>
<intersection>1320.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>720,1320.5,734,1320.5</points>
<connection>
<GID>1022</GID>
<name>IN_1</name></connection>
<intersection>720 8</intersection></hsegment></shape></wire>
<wire>
<ID>1612</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>629.5,1348,685.5,1348</points>
<connection>
<GID>1108</GID>
<name>OUT_3</name></connection>
<intersection>631 7</intersection>
<intersection>685.5 11</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>631,1348,631,1374.5</points>
<intersection>1348 4</intersection>
<intersection>1374.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>631,1374.5,634,1374.5</points>
<connection>
<GID>1270</GID>
<name>IN_3</name></connection>
<intersection>631 7</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>685.5,1321.5,685.5,1348</points>
<intersection>1321.5 12</intersection>
<intersection>1348 4</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>685.5,1321.5,733,1321.5</points>
<intersection>685.5 11</intersection>
<intersection>733 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>733,1314.5,733,1321.5</points>
<intersection>1314.5 14</intersection>
<intersection>1321.5 12</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>733,1314.5,734,1314.5</points>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection>
<intersection>733 13</intersection></hsegment></shape></wire>
<wire>
<ID>1613</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>629.5,1347,631.5,1347</points>
<connection>
<GID>1108</GID>
<name>OUT_2</name></connection>
<intersection>631.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>631.5,1347,631.5,1373.5</points>
<intersection>1347 5</intersection>
<intersection>1373.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>631.5,1373.5,634,1373.5</points>
<connection>
<GID>1270</GID>
<name>IN_2</name></connection>
<intersection>631.5 9</intersection>
<intersection>632 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>632,1373.5,632,1390.5</points>
<intersection>1373.5 10</intersection>
<intersection>1390.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>632,1390.5,634.5,1390.5</points>
<connection>
<GID>1326</GID>
<name>IN_2</name></connection>
<intersection>632 13</intersection></hsegment></shape></wire>
<wire>
<ID>1614</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>629.5,1346,632,1346</points>
<connection>
<GID>1108</GID>
<name>OUT_1</name></connection>
<intersection>632 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>632,1346,632,1372.5</points>
<intersection>1346 2</intersection>
<intersection>1372.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>631.5,1372.5,634,1372.5</points>
<connection>
<GID>1270</GID>
<name>IN_1</name></connection>
<intersection>631.5 8</intersection>
<intersection>632 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>631.5,1372.5,631.5,1389.5</points>
<intersection>1372.5 6</intersection>
<intersection>1389.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>631.5,1389.5,634.5,1389.5</points>
<connection>
<GID>1326</GID>
<name>IN_1</name></connection>
<intersection>631.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1615</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>706.5,1353,707,1353</points>
<connection>
<GID>1314</GID>
<name>IN_0</name></connection>
<intersection>706.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>706.5,1351.5,706.5,1353</points>
<connection>
<GID>1177</GID>
<name>OUT_0</name></connection>
<intersection>1353 0</intersection></vsegment></shape></wire>
<wire>
<ID>1616</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>632.5,1345,632.5,1371.5</points>
<intersection>1345 5</intersection>
<intersection>1371.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>629.5,1345,632.5,1345</points>
<connection>
<GID>1108</GID>
<name>OUT_0</name></connection>
<intersection>632.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>631,1371.5,634,1371.5</points>
<connection>
<GID>1270</GID>
<name>IN_0</name></connection>
<intersection>631 8</intersection>
<intersection>632.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>631,1371.5,631,1388.5</points>
<intersection>1371.5 6</intersection>
<intersection>1388.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>631,1388.5,634.5,1388.5</points>
<connection>
<GID>1326</GID>
<name>IN_0</name></connection>
<intersection>631 8</intersection></hsegment></shape></wire>
<wire>
<ID>1617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572.5,1299.5,572.5,1299.5</points>
<connection>
<GID>1082</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1290</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572.5,1322.5,572.5,1322.5</points>
<connection>
<GID>1083</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1289</GID>
<name>ENABLE_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1620</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>706.5,1350.5,706.5,1351</points>
<connection>
<GID>1177</GID>
<name>OUT_1</name></connection>
<intersection>1351 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>706.5,1351,707,1351</points>
<connection>
<GID>1316</GID>
<name>IN_0</name></connection>
<intersection>706.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1621</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>706.5,1349,706.5,1349.5</points>
<connection>
<GID>1177</GID>
<name>OUT_2</name></connection>
<intersection>1349 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>706.5,1349,707,1349</points>
<connection>
<GID>1327</GID>
<name>IN_0</name></connection>
<intersection>706.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1622</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>706.5,1347,706.5,1348.5</points>
<connection>
<GID>1177</GID>
<name>OUT_3</name></connection>
<intersection>1347 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>706.5,1347,707,1347</points>
<connection>
<GID>1331</GID>
<name>IN_0</name></connection>
<intersection>706.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>1625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>663.5,1360,665,1360</points>
<connection>
<GID>847</GID>
<name>IN_1</name></connection>
<intersection>663.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>663.5,1359.5,663.5,1360</points>
<connection>
<GID>1055</GID>
<name>OUT_2</name></connection>
<intersection>1360 1</intersection></vsegment></shape></wire>
<wire>
<ID>1626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1390.5,580,1390.5</points>
<connection>
<GID>1104</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1389.5,580,1389.5</points>
<connection>
<GID>1104</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1628</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1388.5,580,1388.5</points>
<connection>
<GID>1104</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1387.5,580,1387.5</points>
<connection>
<GID>1104</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1386.5,580,1386.5</points>
<connection>
<GID>1104</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1385.5,580,1385.5</points>
<connection>
<GID>1104</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>550,1392.5,550,1400.5</points>
<connection>
<GID>1102</GID>
<name>count_up</name></connection>
<intersection>1392.5 18</intersection>
<intersection>1400.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>547,1400.5,550,1400.5</points>
<connection>
<GID>1111</GID>
<name>OUT_0</name></connection>
<intersection>548 19</intersection>
<intersection>550 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>549,1392.5,550,1392.5</points>
<connection>
<GID>1102</GID>
<name>count_enable</name></connection>
<intersection>550 0</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>548,1396.5,548,1400.5</points>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection>
<intersection>1400.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>1633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1384.5,580,1384.5</points>
<connection>
<GID>1104</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1383.5,580,1383.5</points>
<connection>
<GID>1104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1107</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1352,615.5,1352</points>
<connection>
<GID>1106</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1422</GID>
<name>IN_7</name></connection>
<intersection>612.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>612.5,1341,612.5,1352</points>
<intersection>1341 10</intersection>
<intersection>1352 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>612.5,1341,616,1341</points>
<connection>
<GID>1405</GID>
<name>IN_7</name></connection>
<intersection>612.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1351,615.5,1351</points>
<connection>
<GID>1106</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1422</GID>
<name>IN_6</name></connection>
<intersection>613 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>613,1340,613,1351</points>
<intersection>1340 7</intersection>
<intersection>1351 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>613,1340,616,1340</points>
<connection>
<GID>1405</GID>
<name>IN_6</name></connection>
<intersection>613 6</intersection></hsegment></shape></wire>
<wire>
<ID>1637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1350,615.5,1350</points>
<connection>
<GID>1106</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1422</GID>
<name>IN_5</name></connection>
<intersection>613.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>613.5,1339,613.5,1350</points>
<intersection>1339 7</intersection>
<intersection>1350 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>613.5,1339,616,1339</points>
<connection>
<GID>1405</GID>
<name>IN_5</name></connection>
<intersection>613.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1349,615.5,1349</points>
<connection>
<GID>1106</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1422</GID>
<name>IN_4</name></connection>
<intersection>614 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>614,1338,614,1349</points>
<intersection>1338 7</intersection>
<intersection>1349 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>614,1338,616,1338</points>
<connection>
<GID>1405</GID>
<name>IN_4</name></connection>
<intersection>614 6</intersection></hsegment></shape></wire>
<wire>
<ID>1639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1348,615.5,1348</points>
<connection>
<GID>1106</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1422</GID>
<name>IN_3</name></connection>
<intersection>614.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>614.5,1337,614.5,1348</points>
<intersection>1337 7</intersection>
<intersection>1348 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>614.5,1337,616,1337</points>
<connection>
<GID>1405</GID>
<name>IN_3</name></connection>
<intersection>614.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1640</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1347,615.5,1347</points>
<connection>
<GID>1106</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1422</GID>
<name>IN_2</name></connection>
<intersection>615 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>615,1336,615,1347</points>
<intersection>1336 7</intersection>
<intersection>1347 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>615,1336,616,1336</points>
<connection>
<GID>1405</GID>
<name>IN_2</name></connection>
<intersection>615 6</intersection></hsegment></shape></wire>
<wire>
<ID>1641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1346,615.5,1346</points>
<connection>
<GID>1106</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1422</GID>
<name>IN_1</name></connection>
<intersection>615.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>615.5,1335,615.5,1346</points>
<intersection>1335 7</intersection>
<intersection>1346 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>615.5,1335,616,1335</points>
<connection>
<GID>1405</GID>
<name>IN_1</name></connection>
<intersection>615.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1642</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>612,1345,616,1345</points>
<connection>
<GID>1106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection>
<intersection>616 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>616,1334,616,1345</points>
<connection>
<GID>1405</GID>
<name>IN_0</name></connection>
<intersection>1345 1</intersection></vsegment></shape></wire>
<wire>
<ID>1644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>550,1362.5,550,1381.5</points>
<connection>
<GID>1102</GID>
<name>clear</name></connection>
<intersection>1362.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>550,1362.5,619.5,1362.5</points>
<intersection>550 0</intersection>
<intersection>554 15</intersection>
<intersection>571.5 3</intersection>
<intersection>602 7</intersection>
<intersection>619.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>571.5,1362.5,571.5,1381.5</points>
<connection>
<GID>1104</GID>
<name>clear</name></connection>
<intersection>1362.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>619.5,1342,619.5,1362.5</points>
<intersection>1342 9</intersection>
<intersection>1362.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>602,1343,602,1362.5</points>
<intersection>1343 10</intersection>
<intersection>1362.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>619.5,1342,626.5,1342</points>
<intersection>619.5 6</intersection>
<intersection>626.5 18</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>602,1343,609,1343</points>
<connection>
<GID>1106</GID>
<name>clear</name></connection>
<intersection>602 7</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>554,1358.5,554,1362.5</points>
<connection>
<GID>1114</GID>
<name>OUT_0</name></connection>
<intersection>1362.5 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>626.5,1342,626.5,1343</points>
<connection>
<GID>1108</GID>
<name>clear</name></connection>
<intersection>1342 9</intersection></vsegment></shape></wire>
<wire>
<ID>1645</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>591,1353.5,591,1387.5</points>
<intersection>1353.5 4</intersection>
<intersection>1387.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>576.5,1353.5,591,1353.5</points>
<connection>
<GID>1126</GID>
<name>ENABLE_0</name></connection>
<intersection>591 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>590,1387.5,597,1387.5</points>
<connection>
<GID>1107</GID>
<name>write_enable</name></connection>
<intersection>591 3</intersection>
<intersection>597 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>597,1385.5,597,1393</points>
<connection>
<GID>1457</GID>
<name>IN_0</name></connection>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection>
<intersection>1387.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>1646</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1346,589.5,1346</points>
<connection>
<GID>1126</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1125</GID>
<name>IN_1</name></connection>
<intersection>587.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>587.5,1346,587.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_1</name></connection>
<intersection>1346 1</intersection></vsegment></shape></wire>
<wire>
<ID>1647</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1347,589.5,1347</points>
<connection>
<GID>1126</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1125</GID>
<name>IN_2</name></connection>
<intersection>586.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>586.5,1347,586.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_2</name></connection>
<intersection>1347 1</intersection></vsegment></shape></wire>
<wire>
<ID>1648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1348,589.5,1348</points>
<connection>
<GID>1126</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1125</GID>
<name>IN_3</name></connection>
<intersection>585.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>585.5,1348,585.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_3</name></connection>
<intersection>1348 1</intersection></vsegment></shape></wire>
<wire>
<ID>1649</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1349,589.5,1349</points>
<connection>
<GID>1126</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1125</GID>
<name>IN_4</name></connection>
<intersection>584.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>584.5,1349,584.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_4</name></connection>
<intersection>1349 1</intersection></vsegment></shape></wire>
<wire>
<ID>1650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1350,589.5,1350</points>
<connection>
<GID>1126</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1125</GID>
<name>IN_5</name></connection>
<intersection>583.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>583.5,1350,583.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_5</name></connection>
<intersection>1350 1</intersection></vsegment></shape></wire>
<wire>
<ID>1651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1351,589.5,1351</points>
<connection>
<GID>1126</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1125</GID>
<name>IN_6</name></connection>
<intersection>582.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>582.5,1351,582.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_6</name></connection>
<intersection>1351 1</intersection></vsegment></shape></wire>
<wire>
<ID>1652</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1352,589.5,1352</points>
<connection>
<GID>1126</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1125</GID>
<name>IN_7</name></connection>
<intersection>581.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>581.5,1352,581.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_7</name></connection>
<intersection>1352 1</intersection></vsegment></shape></wire>
<wire>
<ID>1653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1350,604,1350</points>
<connection>
<GID>1106</GID>
<name>IN_5</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_5</name></connection>
<intersection>596 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>596,1340,596,1350</points>
<intersection>1340 6</intersection>
<intersection>1350 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1340,596,1340</points>
<connection>
<GID>1439</GID>
<name>OUT_5</name></connection>
<intersection>596 5</intersection></hsegment></shape></wire>
<wire>
<ID>1654</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1345,604,1345</points>
<connection>
<GID>1106</GID>
<name>IN_0</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_0</name></connection>
<intersection>601 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>601,1335,601,1345</points>
<intersection>1335 6</intersection>
<intersection>1345 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1335,601,1335</points>
<connection>
<GID>1439</GID>
<name>OUT_0</name></connection>
<intersection>601 5</intersection></hsegment></shape></wire>
<wire>
<ID>1655</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1346,604,1346</points>
<connection>
<GID>1106</GID>
<name>IN_1</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_1</name></connection>
<intersection>600 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>600,1336,600,1346</points>
<intersection>1336 6</intersection>
<intersection>1346 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1336,600,1336</points>
<connection>
<GID>1439</GID>
<name>OUT_1</name></connection>
<intersection>600 5</intersection></hsegment></shape></wire>
<wire>
<ID>1656</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1347,604,1347</points>
<connection>
<GID>1106</GID>
<name>IN_2</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_2</name></connection>
<intersection>599 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>599,1337,599,1347</points>
<intersection>1337 6</intersection>
<intersection>1347 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1337,599,1337</points>
<connection>
<GID>1439</GID>
<name>OUT_2</name></connection>
<intersection>599 5</intersection></hsegment></shape></wire>
<wire>
<ID>1657</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1348,604,1348</points>
<connection>
<GID>1106</GID>
<name>IN_3</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_3</name></connection>
<intersection>598 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>598,1338,598,1348</points>
<intersection>1338 6</intersection>
<intersection>1348 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1338,598,1338</points>
<connection>
<GID>1439</GID>
<name>OUT_3</name></connection>
<intersection>598 5</intersection></hsegment></shape></wire>
<wire>
<ID>1658</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1349,604,1349</points>
<connection>
<GID>1106</GID>
<name>IN_4</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_4</name></connection>
<intersection>597 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>597,1339,597,1349</points>
<intersection>1339 6</intersection>
<intersection>1349 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1339,597,1339</points>
<connection>
<GID>1439</GID>
<name>OUT_4</name></connection>
<intersection>597 5</intersection></hsegment></shape></wire>
<wire>
<ID>1659</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1352,604,1352</points>
<connection>
<GID>1106</GID>
<name>IN_7</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_7</name></connection>
<intersection>594 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>594,1342,594,1352</points>
<intersection>1342 6</intersection>
<intersection>1352 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1342,594,1342</points>
<connection>
<GID>1439</GID>
<name>OUT_7</name></connection>
<intersection>594 5</intersection></hsegment></shape></wire>
<wire>
<ID>1660</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>593.5,1351,604,1351</points>
<connection>
<GID>1106</GID>
<name>IN_6</name></connection>
<connection>
<GID>1125</GID>
<name>OUT_6</name></connection>
<intersection>595 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>595,1341,595,1351</points>
<intersection>1341 6</intersection>
<intersection>1351 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>593.5,1341,595,1341</points>
<connection>
<GID>1439</GID>
<name>OUT_6</name></connection>
<intersection>595 5</intersection></hsegment></shape></wire>
<wire>
<ID>1661</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578.5,1345,589.5,1345</points>
<connection>
<GID>1126</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1125</GID>
<name>IN_0</name></connection>
<intersection>588.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>588.5,1345,588.5,1380</points>
<connection>
<GID>1107</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>1107</GID>
<name>DATA_IN_0</name></connection>
<intersection>1345 1</intersection></vsegment></shape></wire>
<wire>
<ID>1664</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>706.5,1337,707,1337</points>
<connection>
<GID>1332</GID>
<name>IN_0</name></connection>
<intersection>706.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>706.5,1335.5,706.5,1337</points>
<connection>
<GID>1179</GID>
<name>OUT_0</name></connection>
<intersection>1337 1</intersection></vsegment></shape></wire>
<wire>
<ID>1665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571.5,1333,625,1333</points>
<intersection>571.5 8</intersection>
<intersection>625 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>625,1285.5,625,1333</points>
<intersection>1285.5 18</intersection>
<intersection>1290.5 19</intersection>
<intersection>1295.5 20</intersection>
<intersection>1300.5 21</intersection>
<intersection>1305.5 22</intersection>
<intersection>1310.5 23</intersection>
<intersection>1315.5 24</intersection>
<intersection>1320.5 25</intersection>
<intersection>1333 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>571.5,1328.5,571.5,1333</points>
<intersection>1328.5 10</intersection>
<intersection>1330 27</intersection>
<intersection>1333 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>571.5,1328.5,576,1328.5</points>
<connection>
<GID>1207</GID>
<name>IN_0</name></connection>
<intersection>571.5 8</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>625,1285.5,630.5,1285.5</points>
<connection>
<GID>1178</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>625,1290.5,630.5,1290.5</points>
<connection>
<GID>1176</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>625,1295.5,630.5,1295.5</points>
<connection>
<GID>1173</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>625,1300.5,630.5,1300.5</points>
<connection>
<GID>1171</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>625,1305.5,630.5,1305.5</points>
<connection>
<GID>1168</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>625,1310.5,630.5,1310.5</points>
<connection>
<GID>1163</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>625,1315.5,630.5,1315.5</points>
<connection>
<GID>1161</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>625,1320.5,630.5,1320.5</points>
<connection>
<GID>1158</GID>
<name>SEL_0</name></connection>
<intersection>625 7</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>570,1330,571.5,1330</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>571.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>583,1299.5,583,1328.5</points>
<intersection>1299.5 2</intersection>
<intersection>1328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582,1328.5,583,1328.5</points>
<connection>
<GID>1207</GID>
<name>OUT_0</name></connection>
<intersection>583 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>583,1299.5,587.5,1299.5</points>
<connection>
<GID>1134</GID>
<name>ENABLE_0</name></connection>
<intersection>583 0</intersection></hsegment></shape></wire>
<wire>
<ID>1667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>587.5,1322.5,587.5,1329.5</points>
<connection>
<GID>1133</GID>
<name>ENABLE_0</name></connection>
<intersection>1329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>582,1329.5,587.5,1329.5</points>
<connection>
<GID>1207</GID>
<name>OUT_1</name></connection>
<intersection>587.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1668</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>604,1286.5,604,1287</points>
<connection>
<GID>1216</GID>
<name>carry_in</name></connection>
<connection>
<GID>1215</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>1669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597.5,1283,597.5,1300</points>
<intersection>1283 2</intersection>
<intersection>1300 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597.5,1300,601,1300</points>
<connection>
<GID>1215</GID>
<name>IN_B_0</name></connection>
<intersection>597.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1283,597.5,1283</points>
<connection>
<GID>1134</GID>
<name>OUT_0</name></connection>
<intersection>597.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>597,1285,597,1299</points>
<intersection>1285 2</intersection>
<intersection>1299 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>597,1299,601,1299</points>
<connection>
<GID>1215</GID>
<name>IN_B_1</name></connection>
<intersection>597 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1285,597,1285</points>
<connection>
<GID>1134</GID>
<name>OUT_2</name></connection>
<intersection>597 0</intersection></hsegment></shape></wire>
<wire>
<ID>1671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,1287,596.5,1298</points>
<intersection>1287 2</intersection>
<intersection>1298 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596.5,1298,601,1298</points>
<connection>
<GID>1215</GID>
<name>IN_B_2</name></connection>
<intersection>596.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1287,596.5,1287</points>
<connection>
<GID>1134</GID>
<name>OUT_4</name></connection>
<intersection>596.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596,1289,596,1297</points>
<intersection>1289 2</intersection>
<intersection>1297 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596,1297,601,1297</points>
<connection>
<GID>1215</GID>
<name>IN_B_3</name></connection>
<intersection>596 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1289,596,1289</points>
<connection>
<GID>1134</GID>
<name>OUT_6</name></connection>
<intersection>596 0</intersection></hsegment></shape></wire>
<wire>
<ID>1673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593.5,1283.5,593.5,1291</points>
<intersection>1283.5 1</intersection>
<intersection>1291 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>593.5,1283.5,601,1283.5</points>
<connection>
<GID>1216</GID>
<name>IN_B_0</name></connection>
<intersection>593.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1291,593.5,1291</points>
<connection>
<GID>1134</GID>
<name>OUT_8</name></connection>
<intersection>593.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,1282.5,592.5,1293</points>
<intersection>1282.5 1</intersection>
<intersection>1293 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,1282.5,601,1282.5</points>
<connection>
<GID>1216</GID>
<name>IN_B_1</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1293,592.5,1293</points>
<connection>
<GID>1134</GID>
<name>OUT_10</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591.5,1281.5,591.5,1295</points>
<intersection>1281.5 1</intersection>
<intersection>1295 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591.5,1281.5,601,1281.5</points>
<connection>
<GID>1216</GID>
<name>IN_B_2</name></connection>
<intersection>591.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1295,591.5,1295</points>
<connection>
<GID>1134</GID>
<name>OUT_12</name></connection>
<intersection>591.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,1280.5,590.5,1297</points>
<intersection>1280.5 1</intersection>
<intersection>1297 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,1280.5,601,1280.5</points>
<connection>
<GID>1216</GID>
<name>IN_B_3</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1297,590.5,1297</points>
<connection>
<GID>1134</GID>
<name>OUT_14</name></connection>
<intersection>590.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>595.5,1284,595.5,1293</points>
<intersection>1284 2</intersection>
<intersection>1293 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595.5,1293,601,1293</points>
<connection>
<GID>1215</GID>
<name>IN_0</name></connection>
<intersection>595.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1284,595.5,1284</points>
<connection>
<GID>1134</GID>
<name>OUT_1</name></connection>
<intersection>595.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>595,1286,595,1292</points>
<intersection>1286 2</intersection>
<intersection>1292 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595,1292,601,1292</points>
<connection>
<GID>1215</GID>
<name>IN_1</name></connection>
<intersection>595 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1286,595,1286</points>
<connection>
<GID>1134</GID>
<name>OUT_3</name></connection>
<intersection>595 0</intersection></hsegment></shape></wire>
<wire>
<ID>1679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594.5,1288,594.5,1291</points>
<intersection>1288 2</intersection>
<intersection>1291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594.5,1291,601,1291</points>
<connection>
<GID>1215</GID>
<name>IN_2</name></connection>
<intersection>594.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1288,594.5,1288</points>
<connection>
<GID>1134</GID>
<name>OUT_5</name></connection>
<intersection>594.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1680</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>589.5,1290,601,1290</points>
<connection>
<GID>1134</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1215</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,1276.5,593,1292</points>
<intersection>1276.5 1</intersection>
<intersection>1292 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>593,1276.5,601,1276.5</points>
<connection>
<GID>1216</GID>
<name>IN_0</name></connection>
<intersection>593 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1292,593,1292</points>
<connection>
<GID>1134</GID>
<name>OUT_9</name></connection>
<intersection>593 0</intersection></hsegment></shape></wire>
<wire>
<ID>1682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592,1275.5,592,1294</points>
<intersection>1275.5 1</intersection>
<intersection>1294 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592,1275.5,601,1275.5</points>
<connection>
<GID>1216</GID>
<name>IN_1</name></connection>
<intersection>592 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1294,592,1294</points>
<connection>
<GID>1134</GID>
<name>OUT_11</name></connection>
<intersection>592 0</intersection></hsegment></shape></wire>
<wire>
<ID>1683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591,1274.5,591,1296</points>
<intersection>1274.5 1</intersection>
<intersection>1296 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591,1274.5,601,1274.5</points>
<connection>
<GID>1216</GID>
<name>IN_2</name></connection>
<intersection>591 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1296,591,1296</points>
<connection>
<GID>1134</GID>
<name>OUT_13</name></connection>
<intersection>591 0</intersection></hsegment></shape></wire>
<wire>
<ID>1684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,1273.5,590,1298</points>
<intersection>1273.5 1</intersection>
<intersection>1298 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,1273.5,601,1273.5</points>
<connection>
<GID>1216</GID>
<name>IN_3</name></connection>
<intersection>590 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1298,590,1298</points>
<connection>
<GID>1134</GID>
<name>OUT_15</name></connection>
<intersection>590 0</intersection></hsegment></shape></wire>
<wire>
<ID>1685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594.5,1304,594.5,1306</points>
<intersection>1304 1</intersection>
<intersection>1306 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594.5,1304,597.5,1304</points>
<connection>
<GID>1185</GID>
<name>IN_1</name></connection>
<intersection>594.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1306,594.5,1306</points>
<connection>
<GID>1133</GID>
<name>OUT_0</name></connection>
<intersection>594.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1686</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>595,1306,597.5,1306</points>
<connection>
<GID>1185</GID>
<name>IN_0</name></connection>
<intersection>595 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>595,1306,595,1307</points>
<intersection>1306 1</intersection>
<intersection>1307 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>589.5,1307,595,1307</points>
<connection>
<GID>1133</GID>
<name>OUT_1</name></connection>
<intersection>595 3</intersection></hsegment></shape></wire>
<wire>
<ID>1687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>595.5,1307.5,595.5,1308</points>
<intersection>1307.5 1</intersection>
<intersection>1308 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>595.5,1307.5,602.5,1307.5</points>
<connection>
<GID>1196</GID>
<name>IN_1</name></connection>
<intersection>595.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1308,595.5,1308</points>
<connection>
<GID>1133</GID>
<name>OUT_2</name></connection>
<intersection>595.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1688</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>595.5,1309.5,602.5,1309.5</points>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection>
<intersection>595.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>595.5,1309,595.5,1309.5</points>
<intersection>1309 4</intersection>
<intersection>1309.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>589.5,1309,595.5,1309</points>
<connection>
<GID>1133</GID>
<name>OUT_3</name></connection>
<intersection>595.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1689</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>589.5,1310,595,1310</points>
<connection>
<GID>1133</GID>
<name>OUT_4</name></connection>
<intersection>595 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>595,1310,595,1311</points>
<intersection>1310 1</intersection>
<intersection>1311 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>595,1311,597.5,1311</points>
<connection>
<GID>1211</GID>
<name>IN_1</name></connection>
<intersection>595 5</intersection></hsegment></shape></wire>
<wire>
<ID>1690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594.5,1311,594.5,1313</points>
<intersection>1311 2</intersection>
<intersection>1313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594.5,1313,597.5,1313</points>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection>
<intersection>594.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1311,594.5,1311</points>
<connection>
<GID>1133</GID>
<name>OUT_5</name></connection>
<intersection>594.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594,1312,594,1314.5</points>
<intersection>1312 2</intersection>
<intersection>1314.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>594,1314.5,602.5,1314.5</points>
<connection>
<GID>1225</GID>
<name>IN_1</name></connection>
<intersection>594 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1312,594,1312</points>
<connection>
<GID>1133</GID>
<name>OUT_6</name></connection>
<intersection>594 0</intersection></hsegment></shape></wire>
<wire>
<ID>1692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593.5,1313,593.5,1316.5</points>
<intersection>1313 2</intersection>
<intersection>1316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>593.5,1316.5,602.5,1316.5</points>
<connection>
<GID>1225</GID>
<name>IN_0</name></connection>
<intersection>593.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1313,593.5,1313</points>
<connection>
<GID>1133</GID>
<name>OUT_7</name></connection>
<intersection>593.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,1314,593,1318</points>
<intersection>1314 2</intersection>
<intersection>1318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>593,1318,597.5,1318</points>
<connection>
<GID>1234</GID>
<name>IN_1</name></connection>
<intersection>593 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1314,593,1314</points>
<connection>
<GID>1133</GID>
<name>OUT_8</name></connection>
<intersection>593 0</intersection></hsegment></shape></wire>
<wire>
<ID>1694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,1315,592.5,1320</points>
<intersection>1315 2</intersection>
<intersection>1320 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,1320,597.5,1320</points>
<connection>
<GID>1234</GID>
<name>IN_0</name></connection>
<intersection>592.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1315,592.5,1315</points>
<connection>
<GID>1133</GID>
<name>OUT_9</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592,1316,592,1321.5</points>
<intersection>1316 2</intersection>
<intersection>1321.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592,1321.5,602.5,1321.5</points>
<connection>
<GID>1095</GID>
<name>IN_1</name></connection>
<intersection>592 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1316,592,1316</points>
<connection>
<GID>1133</GID>
<name>OUT_10</name></connection>
<intersection>592 0</intersection></hsegment></shape></wire>
<wire>
<ID>1696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591.5,1317,591.5,1323.5</points>
<intersection>1317 2</intersection>
<intersection>1323.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591.5,1323.5,602.5,1323.5</points>
<connection>
<GID>1095</GID>
<name>IN_0</name></connection>
<intersection>591.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1317,591.5,1317</points>
<connection>
<GID>1133</GID>
<name>OUT_11</name></connection>
<intersection>591.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591,1318,591,1325</points>
<intersection>1318 2</intersection>
<intersection>1325 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>591,1325,597.5,1325</points>
<connection>
<GID>1098</GID>
<name>IN_1</name></connection>
<intersection>591 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1318,591,1318</points>
<connection>
<GID>1133</GID>
<name>OUT_12</name></connection>
<intersection>591 0</intersection></hsegment></shape></wire>
<wire>
<ID>1698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590.5,1319,590.5,1327</points>
<intersection>1319 2</intersection>
<intersection>1327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590.5,1327,597.5,1327</points>
<connection>
<GID>1098</GID>
<name>IN_0</name></connection>
<intersection>590.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1319,590.5,1319</points>
<connection>
<GID>1133</GID>
<name>OUT_13</name></connection>
<intersection>590.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,1320,590,1328.5</points>
<intersection>1320 2</intersection>
<intersection>1328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,1328.5,602.5,1328.5</points>
<connection>
<GID>1101</GID>
<name>IN_1</name></connection>
<intersection>590 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>589.5,1320,590,1320</points>
<connection>
<GID>1133</GID>
<name>OUT_14</name></connection>
<intersection>590 0</intersection></hsegment></shape></wire>
<wire>
<ID>1700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>589.5,1321,589.5,1330.5</points>
<connection>
<GID>1133</GID>
<name>OUT_15</name></connection>
<intersection>1330.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589.5,1330.5,602.5,1330.5</points>
<connection>
<GID>1101</GID>
<name>IN_0</name></connection>
<intersection>589.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1282,618.5,1296.5</points>
<intersection>1282 1</intersection>
<intersection>1296.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1282,628.5,1282</points>
<connection>
<GID>1178</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1296.5,618.5,1296.5</points>
<connection>
<GID>1215</GID>
<name>OUT_0</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1287,618.5,1295.5</points>
<intersection>1287 1</intersection>
<intersection>1295.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1287,628.5,1287</points>
<connection>
<GID>1176</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1295.5,618.5,1295.5</points>
<connection>
<GID>1215</GID>
<name>OUT_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1292,618.5,1294.5</points>
<intersection>1292 1</intersection>
<intersection>1294.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1292,628.5,1292</points>
<connection>
<GID>1173</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1294.5,618.5,1294.5</points>
<connection>
<GID>1215</GID>
<name>OUT_2</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1293.5,618.5,1297</points>
<intersection>1293.5 2</intersection>
<intersection>1297 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1297,628.5,1297</points>
<connection>
<GID>1171</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1293.5,618.5,1293.5</points>
<connection>
<GID>1215</GID>
<name>OUT_3</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1280,618.5,1302</points>
<intersection>1280 2</intersection>
<intersection>1302 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1302,628.5,1302</points>
<connection>
<GID>1168</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1280,618.5,1280</points>
<connection>
<GID>1216</GID>
<name>OUT_0</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1279,618.5,1307</points>
<intersection>1279 2</intersection>
<intersection>1307 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1307,628.5,1307</points>
<connection>
<GID>1163</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1279,618.5,1279</points>
<connection>
<GID>1216</GID>
<name>OUT_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1278,618.5,1312</points>
<intersection>1278 2</intersection>
<intersection>1312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1312,628.5,1312</points>
<connection>
<GID>1161</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1278,618.5,1278</points>
<connection>
<GID>1216</GID>
<name>OUT_2</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1708</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1277,618.5,1317</points>
<intersection>1277 2</intersection>
<intersection>1317 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,1317,628.5,1317</points>
<connection>
<GID>1158</GID>
<name>IN_0</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>609,1277,618.5,1277</points>
<connection>
<GID>1216</GID>
<name>OUT_3</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,1284,616,1305</points>
<intersection>1284 1</intersection>
<intersection>1305 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616,1284,628.5,1284</points>
<connection>
<GID>1178</GID>
<name>IN_1</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>603.5,1305,616,1305</points>
<connection>
<GID>1185</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>1710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1289,618.5,1308.5</points>
<intersection>1289 2</intersection>
<intersection>1308.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608.5,1308.5,618.5,1308.5</points>
<connection>
<GID>1196</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>618.5,1289,628.5,1289</points>
<connection>
<GID>1176</GID>
<name>IN_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,1294,616,1312</points>
<intersection>1294 2</intersection>
<intersection>1312 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603.5,1312,616,1312</points>
<connection>
<GID>1211</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>616,1294,628.5,1294</points>
<connection>
<GID>1173</GID>
<name>IN_1</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>1712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1299,618.5,1315.5</points>
<intersection>1299 2</intersection>
<intersection>1315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608.5,1315.5,618.5,1315.5</points>
<connection>
<GID>1225</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>618.5,1299,628.5,1299</points>
<connection>
<GID>1171</GID>
<name>IN_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,1304,616,1319</points>
<intersection>1304 2</intersection>
<intersection>1319 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603.5,1319,616,1319</points>
<connection>
<GID>1234</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>616,1304,628.5,1304</points>
<connection>
<GID>1168</GID>
<name>IN_1</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>1714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1309,618.5,1322.5</points>
<intersection>1309 2</intersection>
<intersection>1322.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608.5,1322.5,618.5,1322.5</points>
<connection>
<GID>1095</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>618.5,1309,628.5,1309</points>
<connection>
<GID>1163</GID>
<name>IN_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,1314,616,1326</points>
<intersection>1314 2</intersection>
<intersection>1326 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>603.5,1326,616,1326</points>
<connection>
<GID>1098</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>616,1314,628.5,1314</points>
<connection>
<GID>1161</GID>
<name>IN_1</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>1716</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,1319,618.5,1329.5</points>
<intersection>1319 2</intersection>
<intersection>1329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>608.5,1329.5,618.5,1329.5</points>
<connection>
<GID>1101</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>618.5,1319,628.5,1319</points>
<connection>
<GID>1158</GID>
<name>IN_1</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1283,640,1296.5</points>
<intersection>1283 2</intersection>
<intersection>1296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1296.5,671.5,1296.5</points>
<connection>
<GID>1180</GID>
<name>IN_0</name></connection>
<intersection>640 0</intersection>
<intersection>641 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1283,640,1283</points>
<connection>
<GID>1178</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>641,1292.5,641,1296.5</points>
<intersection>1292.5 8</intersection>
<intersection>1296.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>641,1292.5,662,1292.5</points>
<intersection>641 7</intersection>
<intersection>662 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>662,1276,662,1292.5</points>
<connection>
<GID>1202</GID>
<name>N_in2</name></connection>
<intersection>1276 13</intersection>
<intersection>1292.5 8</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>662,1276,669.5,1276</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>662 9</intersection></hsegment></shape></wire>
<wire>
<ID>1718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1288,640,1297.5</points>
<intersection>1288 2</intersection>
<intersection>1297.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1297.5,671.5,1297.5</points>
<connection>
<GID>1180</GID>
<name>IN_1</name></connection>
<intersection>640 0</intersection>
<intersection>641.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1288,640,1288</points>
<connection>
<GID>1176</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>641.5,1293,641.5,1297.5</points>
<intersection>1293 8</intersection>
<intersection>1297.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>641.5,1293,659.5,1293</points>
<intersection>641.5 7</intersection>
<intersection>659.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>659.5,1277,659.5,1293</points>
<connection>
<GID>1200</GID>
<name>N_in2</name></connection>
<intersection>1277 15</intersection>
<intersection>1293 8</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>659.5,1277,669.5,1277</points>
<connection>
<GID>1513</GID>
<name>IN_1</name></connection>
<intersection>659.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>1719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1293,640,1298.5</points>
<intersection>1293 2</intersection>
<intersection>1298.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1298.5,671.5,1298.5</points>
<connection>
<GID>1180</GID>
<name>IN_2</name></connection>
<intersection>640 0</intersection>
<intersection>642 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1293,640,1293</points>
<connection>
<GID>1173</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>642,1293.5,642,1298.5</points>
<intersection>1293.5 8</intersection>
<intersection>1298.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>642,1293.5,657,1293.5</points>
<intersection>642 7</intersection>
<intersection>657 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>657,1278,657,1293.5</points>
<connection>
<GID>1198</GID>
<name>N_in2</name></connection>
<intersection>1278 15</intersection>
<intersection>1293.5 8</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>657,1278,669.5,1278</points>
<connection>
<GID>1513</GID>
<name>IN_2</name></connection>
<intersection>657 9</intersection></hsegment></shape></wire>
<wire>
<ID>1720</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,1299.5,671.5,1299.5</points>
<connection>
<GID>1180</GID>
<name>IN_3</name></connection>
<intersection>640 20</intersection>
<intersection>642.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>642.5,1294,642.5,1299.5</points>
<intersection>1294 9</intersection>
<intersection>1299.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>642.5,1294,654.5,1294</points>
<intersection>642.5 8</intersection>
<intersection>654.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>654.5,1279,654.5,1294</points>
<connection>
<GID>1195</GID>
<name>N_in2</name></connection>
<intersection>1279 16</intersection>
<intersection>1294 9</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>654.5,1279,669.5,1279</points>
<connection>
<GID>1513</GID>
<name>IN_3</name></connection>
<intersection>654.5 10</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>640,1298,640,1299.5</points>
<intersection>1298 21</intersection>
<intersection>1299.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>632.5,1298,640,1298</points>
<connection>
<GID>1171</GID>
<name>OUT</name></connection>
<intersection>640 20</intersection></hsegment></shape></wire>
<wire>
<ID>1721</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1300.5,640,1303</points>
<intersection>1300.5 1</intersection>
<intersection>1303 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1300.5,671.5,1300.5</points>
<connection>
<GID>1180</GID>
<name>IN_4</name></connection>
<intersection>640 0</intersection>
<intersection>643 8</intersection>
<intersection>668 15</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1303,640,1303</points>
<connection>
<GID>1168</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>643,1294.5,643,1300.5</points>
<intersection>1294.5 9</intersection>
<intersection>1300.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>643,1294.5,652,1294.5</points>
<intersection>643 8</intersection>
<intersection>652 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>652,1292,652,1294.5</points>
<connection>
<GID>1193</GID>
<name>N_in2</name></connection>
<intersection>1294.5 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>668,1280,668,1300.5</points>
<intersection>1280 16</intersection>
<intersection>1300.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>668,1280,669.5,1280</points>
<connection>
<GID>1513</GID>
<name>IN_4</name></connection>
<intersection>668 15</intersection></hsegment></shape></wire>
<wire>
<ID>1722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1301.5,640,1308</points>
<intersection>1301.5 1</intersection>
<intersection>1308 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1301.5,671.5,1301.5</points>
<connection>
<GID>1180</GID>
<name>IN_5</name></connection>
<intersection>640 0</intersection>
<intersection>643.5 7</intersection>
<intersection>668.5 14</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1308,640,1308</points>
<connection>
<GID>1163</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>643.5,1295,643.5,1301.5</points>
<intersection>1295 8</intersection>
<intersection>1301.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>643.5,1295,649.5,1295</points>
<intersection>643.5 7</intersection>
<intersection>649.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>649.5,1292,649.5,1295</points>
<connection>
<GID>1191</GID>
<name>N_in2</name></connection>
<intersection>1295 8</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>668.5,1281,668.5,1301.5</points>
<intersection>1281 15</intersection>
<intersection>1301.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>668.5,1281,669.5,1281</points>
<connection>
<GID>1513</GID>
<name>IN_5</name></connection>
<intersection>668.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>1723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1302.5,640,1313</points>
<intersection>1302.5 1</intersection>
<intersection>1313 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>640,1302.5,671.5,1302.5</points>
<connection>
<GID>1180</GID>
<name>IN_6</name></connection>
<intersection>640 0</intersection>
<intersection>644 7</intersection>
<intersection>669 14</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1313,640,1313</points>
<connection>
<GID>1161</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>644,1295.5,644,1302.5</points>
<intersection>1295.5 8</intersection>
<intersection>1302.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>644,1295.5,647,1295.5</points>
<intersection>644 7</intersection>
<intersection>647 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>647,1292,647,1295.5</points>
<connection>
<GID>1189</GID>
<name>N_in2</name></connection>
<intersection>1295.5 8</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>669,1282,669,1302.5</points>
<intersection>1282 15</intersection>
<intersection>1302.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>669,1282,669.5,1282</points>
<connection>
<GID>1513</GID>
<name>IN_6</name></connection>
<intersection>669 14</intersection></hsegment></shape></wire>
<wire>
<ID>1724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>640,1303.5,640,1318</points>
<intersection>1303.5 2</intersection>
<intersection>1318 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>632.5,1318,640,1318</points>
<connection>
<GID>1158</GID>
<name>OUT</name></connection>
<intersection>640 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>640,1303.5,671.5,1303.5</points>
<connection>
<GID>1180</GID>
<name>IN_7</name></connection>
<intersection>640 0</intersection>
<intersection>644.5 5</intersection>
<intersection>669.5 13</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>644.5,1292,644.5,1303.5</points>
<connection>
<GID>1187</GID>
<name>N_in2</name></connection>
<intersection>1303.5 2</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>669.5,1283,669.5,1303.5</points>
<connection>
<GID>1513</GID>
<name>IN_7</name></connection>
<intersection>1303.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1725</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454,1290.5,485,1290.5</points>
<connection>
<GID>1103</GID>
<name>OUT_6</name></connection>
<intersection>472.5 4</intersection>
<intersection>485 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>485,1290.5,485,1330</points>
<connection>
<GID>1160</GID>
<name>IN_3</name></connection>
<intersection>1290.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>472.5,1290.5,472.5,1330</points>
<connection>
<GID>1141</GID>
<name>IN_3</name></connection>
<intersection>1290.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455.5,1319,485,1319</points>
<connection>
<GID>1162</GID>
<name>IN_3</name></connection>
<connection>
<GID>1142</GID>
<name>IN_3</name></connection>
<intersection>455.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>455.5,1289.5,455.5,1319</points>
<intersection>1289.5 5</intersection>
<intersection>1319 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1289.5,455.5,1289.5</points>
<connection>
<GID>1103</GID>
<name>OUT_5</name></connection>
<intersection>455.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1727</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456,1309.5,485,1309.5</points>
<connection>
<GID>1164</GID>
<name>IN_3</name></connection>
<connection>
<GID>1143</GID>
<name>IN_3</name></connection>
<intersection>456 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>456,1288.5,456,1309.5</points>
<intersection>1288.5 6</intersection>
<intersection>1309.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>454,1288.5,456,1288.5</points>
<connection>
<GID>1103</GID>
<name>OUT_4</name></connection>
<intersection>456 4</intersection></hsegment></shape></wire>
<wire>
<ID>1728</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456.5,1298.5,485,1298.5</points>
<connection>
<GID>1165</GID>
<name>IN_3</name></connection>
<connection>
<GID>1144</GID>
<name>IN_3</name></connection>
<intersection>456.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>456.5,1287.5,456.5,1298.5</points>
<intersection>1287.5 5</intersection>
<intersection>1298.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1287.5,456.5,1287.5</points>
<connection>
<GID>1103</GID>
<name>OUT_3</name></connection>
<intersection>456.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1729</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>457.5,1277,485,1277</points>
<connection>
<GID>1146</GID>
<name>IN_3</name></connection>
<connection>
<GID>1167</GID>
<name>IN_3</name></connection>
<intersection>457.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>457.5,1277,457.5,1285.5</points>
<intersection>1277 1</intersection>
<intersection>1285.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1285.5,457.5,1285.5</points>
<connection>
<GID>1103</GID>
<name>OUT_1</name></connection>
<intersection>457.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1730</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>458,1266,485,1266</points>
<connection>
<GID>1147</GID>
<name>IN_3</name></connection>
<connection>
<GID>1170</GID>
<name>IN_3</name></connection>
<intersection>458 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>458,1266,458,1284.5</points>
<intersection>1266 2</intersection>
<intersection>1284.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1284.5,458,1284.5</points>
<connection>
<GID>1103</GID>
<name>OUT_0</name></connection>
<intersection>458 4</intersection></hsegment></shape></wire>
<wire>
<ID>1731</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>458.5,1339,485,1339</points>
<connection>
<GID>1157</GID>
<name>IN_2</name></connection>
<connection>
<GID>1139</GID>
<name>IN_2</name></connection>
<intersection>458.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>458.5,1304.5,458.5,1339</points>
<intersection>1304.5 5</intersection>
<intersection>1339 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1304.5,458.5,1304.5</points>
<connection>
<GID>1105</GID>
<name>OUT_7</name></connection>
<intersection>458.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1732</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>459,1328,485,1328</points>
<connection>
<GID>1160</GID>
<name>IN_2</name></connection>
<connection>
<GID>1141</GID>
<name>IN_2</name></connection>
<intersection>459 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>459,1303.5,459,1328</points>
<intersection>1303.5 5</intersection>
<intersection>1328 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1303.5,459,1303.5</points>
<connection>
<GID>1105</GID>
<name>OUT_6</name></connection>
<intersection>459 4</intersection></hsegment></shape></wire>
<wire>
<ID>1733</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>459.5,1317,485,1317</points>
<connection>
<GID>1162</GID>
<name>IN_2</name></connection>
<connection>
<GID>1142</GID>
<name>IN_2</name></connection>
<intersection>459.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>459.5,1302.5,459.5,1317</points>
<intersection>1302.5 7</intersection>
<intersection>1317 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>454,1302.5,459.5,1302.5</points>
<connection>
<GID>1105</GID>
<name>OUT_5</name></connection>
<intersection>459.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460,1307.5,485,1307.5</points>
<connection>
<GID>1164</GID>
<name>IN_2</name></connection>
<connection>
<GID>1143</GID>
<name>IN_2</name></connection>
<intersection>460 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>460,1301.5,460,1307.5</points>
<intersection>1301.5 5</intersection>
<intersection>1307.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1301.5,460,1301.5</points>
<connection>
<GID>1105</GID>
<name>OUT_4</name></connection>
<intersection>460 4</intersection></hsegment></shape></wire>
<wire>
<ID>1735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>460.5,1296.5,485,1296.5</points>
<connection>
<GID>1165</GID>
<name>IN_2</name></connection>
<connection>
<GID>1144</GID>
<name>IN_2</name></connection>
<intersection>460.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>460.5,1296.5,460.5,1300.5</points>
<intersection>1296.5 1</intersection>
<intersection>1300.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1300.5,460.5,1300.5</points>
<connection>
<GID>1105</GID>
<name>OUT_3</name></connection>
<intersection>460.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1736</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>461,1285.5,485,1285.5</points>
<connection>
<GID>1166</GID>
<name>IN_2</name></connection>
<connection>
<GID>1145</GID>
<name>IN_2</name></connection>
<intersection>461 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>461,1285.5,461,1299.5</points>
<intersection>1285.5 1</intersection>
<intersection>1299.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1299.5,461,1299.5</points>
<connection>
<GID>1105</GID>
<name>OUT_2</name></connection>
<intersection>461 4</intersection></hsegment></shape></wire>
<wire>
<ID>1737</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>461.5,1275,485,1275</points>
<connection>
<GID>1146</GID>
<name>IN_2</name></connection>
<connection>
<GID>1167</GID>
<name>IN_2</name></connection>
<intersection>461.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>461.5,1275,461.5,1298.5</points>
<intersection>1275 2</intersection>
<intersection>1298.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1298.5,461.5,1298.5</points>
<connection>
<GID>1105</GID>
<name>OUT_1</name></connection>
<intersection>461.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462,1264,485,1264</points>
<connection>
<GID>1147</GID>
<name>IN_2</name></connection>
<connection>
<GID>1170</GID>
<name>IN_2</name></connection>
<intersection>462 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462,1264,462,1297.5</points>
<intersection>1264 1</intersection>
<intersection>1297.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1297.5,462,1297.5</points>
<connection>
<GID>1105</GID>
<name>OUT_0</name></connection>
<intersection>462 4</intersection></hsegment></shape></wire>
<wire>
<ID>1739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462.5,1337,485,1337</points>
<connection>
<GID>1157</GID>
<name>IN_1</name></connection>
<connection>
<GID>1139</GID>
<name>IN_1</name></connection>
<intersection>462.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462.5,1318,462.5,1337</points>
<intersection>1318 5</intersection>
<intersection>1337 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1318,462.5,1318</points>
<connection>
<GID>1136</GID>
<name>OUT_7</name></connection>
<intersection>462.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1740</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>463,1326,485,1326</points>
<connection>
<GID>1160</GID>
<name>IN_1</name></connection>
<connection>
<GID>1141</GID>
<name>IN_1</name></connection>
<intersection>463 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>463,1317,463,1326</points>
<intersection>1317 5</intersection>
<intersection>1326 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1317,463,1317</points>
<connection>
<GID>1136</GID>
<name>OUT_6</name></connection>
<intersection>463 4</intersection></hsegment></shape></wire>
<wire>
<ID>1741</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454,1316,485,1316</points>
<connection>
<GID>1136</GID>
<name>OUT_5</name></connection>
<intersection>472.5 9</intersection>
<intersection>485 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>485,1315,485,1316</points>
<connection>
<GID>1162</GID>
<name>IN_1</name></connection>
<intersection>1316 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>472.5,1315,472.5,1316</points>
<connection>
<GID>1142</GID>
<name>IN_1</name></connection>
<intersection>1316 1</intersection></vsegment></shape></wire>
<wire>
<ID>1742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464,1305.5,485,1305.5</points>
<connection>
<GID>1164</GID>
<name>IN_1</name></connection>
<connection>
<GID>1143</GID>
<name>IN_1</name></connection>
<intersection>464 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>464,1305.5,464,1315</points>
<intersection>1305.5 1</intersection>
<intersection>1315 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1315,464,1315</points>
<connection>
<GID>1136</GID>
<name>OUT_4</name></connection>
<intersection>464 4</intersection></hsegment></shape></wire>
<wire>
<ID>1743</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464.5,1294.5,485,1294.5</points>
<connection>
<GID>1165</GID>
<name>IN_1</name></connection>
<connection>
<GID>1144</GID>
<name>IN_1</name></connection>
<intersection>464.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>464.5,1294.5,464.5,1314</points>
<intersection>1294.5 1</intersection>
<intersection>1314 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1314,464.5,1314</points>
<connection>
<GID>1136</GID>
<name>OUT_3</name></connection>
<intersection>464.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>465,1283.5,485,1283.5</points>
<connection>
<GID>1166</GID>
<name>IN_1</name></connection>
<connection>
<GID>1145</GID>
<name>IN_1</name></connection>
<intersection>465 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>465,1283.5,465,1313</points>
<intersection>1283.5 1</intersection>
<intersection>1313 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1313,465,1313</points>
<connection>
<GID>1136</GID>
<name>OUT_2</name></connection>
<intersection>465 4</intersection></hsegment></shape></wire>
<wire>
<ID>1745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>465.5,1273,485,1273</points>
<connection>
<GID>1146</GID>
<name>IN_1</name></connection>
<connection>
<GID>1167</GID>
<name>IN_1</name></connection>
<intersection>465.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>465.5,1273,465.5,1312</points>
<intersection>1273 1</intersection>
<intersection>1312 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1312,465.5,1312</points>
<connection>
<GID>1136</GID>
<name>OUT_1</name></connection>
<intersection>465.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1746</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>466,1262,485,1262</points>
<connection>
<GID>1147</GID>
<name>IN_1</name></connection>
<connection>
<GID>1170</GID>
<name>IN_1</name></connection>
<intersection>466 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>466,1262,466,1311</points>
<intersection>1262 2</intersection>
<intersection>1311 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1311,466,1311</points>
<connection>
<GID>1136</GID>
<name>OUT_0</name></connection>
<intersection>466 4</intersection></hsegment></shape></wire>
<wire>
<ID>1747</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>466.5,1331,466.5,1335</points>
<intersection>1331 9</intersection>
<intersection>1335 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>466.5,1335,485,1335</points>
<connection>
<GID>1157</GID>
<name>IN_0</name></connection>
<connection>
<GID>1139</GID>
<name>IN_0</name></connection>
<intersection>466.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>454,1331,466.5,1331</points>
<connection>
<GID>1138</GID>
<name>OUT_7</name></connection>
<intersection>466.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1748</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>467,1324,467,1330</points>
<intersection>1324 11</intersection>
<intersection>1330 12</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>467,1324,485,1324</points>
<connection>
<GID>1160</GID>
<name>IN_0</name></connection>
<connection>
<GID>1141</GID>
<name>IN_0</name></connection>
<intersection>467 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>454,1330,467,1330</points>
<connection>
<GID>1138</GID>
<name>OUT_6</name></connection>
<intersection>467 7</intersection></hsegment></shape></wire>
<wire>
<ID>1749</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>467.5,1313,467.5,1329</points>
<intersection>1313 10</intersection>
<intersection>1329 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>467.5,1313,485,1313</points>
<connection>
<GID>1162</GID>
<name>IN_0</name></connection>
<connection>
<GID>1142</GID>
<name>IN_0</name></connection>
<intersection>467.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>454,1329,467.5,1329</points>
<connection>
<GID>1138</GID>
<name>OUT_5</name></connection>
<intersection>467.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1750</ID>
<shape>
<vsegment>
<ID>13</ID>
<points>468,1303.5,468,1328</points>
<intersection>1303.5 16</intersection>
<intersection>1328 17</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>468,1303.5,485,1303.5</points>
<connection>
<GID>1164</GID>
<name>IN_0</name></connection>
<connection>
<GID>1143</GID>
<name>IN_0</name></connection>
<intersection>468 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>454,1328,468,1328</points>
<connection>
<GID>1138</GID>
<name>OUT_4</name></connection>
<intersection>468 13</intersection></hsegment></shape></wire>
<wire>
<ID>1751</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>469,1281.5,469,1326</points>
<intersection>1281.5 7</intersection>
<intersection>1326 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>469,1281.5,485,1281.5</points>
<connection>
<GID>1166</GID>
<name>IN_0</name></connection>
<connection>
<GID>1145</GID>
<name>IN_0</name></connection>
<intersection>469 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>454,1326,469,1326</points>
<connection>
<GID>1138</GID>
<name>OUT_2</name></connection>
<intersection>469 4</intersection></hsegment></shape></wire>
<wire>
<ID>1752</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>469.5,1271,469.5,1325</points>
<intersection>1271 10</intersection>
<intersection>1325 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>469.5,1271,485,1271</points>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection>
<connection>
<GID>1167</GID>
<name>IN_0</name></connection>
<intersection>469.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>454,1325,469.5,1325</points>
<connection>
<GID>1138</GID>
<name>OUT_1</name></connection>
<intersection>469.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1308.5,497,1338</points>
<intersection>1308.5 2</intersection>
<intersection>1317 3</intersection>
<intersection>1338 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,1338,497,1338</points>
<connection>
<GID>1139</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1308.5,509,1308.5</points>
<connection>
<GID>1148</GID>
<name>IN_7</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>497,1317,530,1317</points>
<connection>
<GID>1192</GID>
<name>IN_7</name></connection>
<intersection>497 0</intersection>
<intersection>502 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>502,1317,502,1330</points>
<intersection>1317 3</intersection>
<intersection>1330 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>502,1330,507,1330</points>
<connection>
<GID>1420</GID>
<name>IN_7</name></connection>
<intersection>502 6</intersection></hsegment></shape></wire>
<wire>
<ID>1754</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1307.5,497,1327</points>
<intersection>1307.5 2</intersection>
<intersection>1316 4</intersection>
<intersection>1327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,1327,497,1327</points>
<connection>
<GID>1141</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1307.5,509,1307.5</points>
<connection>
<GID>1148</GID>
<name>IN_6</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>497,1316,530,1316</points>
<connection>
<GID>1192</GID>
<name>IN_6</name></connection>
<intersection>497 0</intersection>
<intersection>502.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>502.5,1316,502.5,1329</points>
<intersection>1316 4</intersection>
<intersection>1329 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>502.5,1329,507,1329</points>
<connection>
<GID>1420</GID>
<name>IN_6</name></connection>
<intersection>502.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1306.5,497,1328</points>
<intersection>1306.5 2</intersection>
<intersection>1315 5</intersection>
<intersection>1328 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>485,1328,507,1328</points>
<connection>
<GID>1420</GID>
<name>IN_5</name></connection>
<intersection>485 8</intersection>
<intersection>497 0</intersection>
<intersection>503 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1306.5,509,1306.5</points>
<connection>
<GID>1148</GID>
<name>IN_5</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>497,1315,530,1315</points>
<connection>
<GID>1192</GID>
<name>IN_5</name></connection>
<intersection>497 0</intersection>
<intersection>503 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>503,1315,503,1328</points>
<intersection>1315 5</intersection>
<intersection>1328 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>485,1316,485,1328</points>
<intersection>1316 9</intersection>
<intersection>1328 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>478.5,1316,485,1316</points>
<connection>
<GID>1142</GID>
<name>OUT</name></connection>
<intersection>485 8</intersection></hsegment></shape></wire>
<wire>
<ID>1756</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>491.5,1305.5,509,1305.5</points>
<connection>
<GID>1148</GID>
<name>IN_4</name></connection>
<intersection>491.5 10</intersection>
<intersection>498 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>498,1305.5,498,1314</points>
<intersection>1305.5 1</intersection>
<intersection>1314 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>498,1314,530,1314</points>
<connection>
<GID>1192</GID>
<name>IN_4</name></connection>
<intersection>498 4</intersection>
<intersection>503.5 11</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>491.5,1305.5,491.5,1306.5</points>
<intersection>1305.5 1</intersection>
<intersection>1306.5 13</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>503.5,1314,503.5,1327</points>
<intersection>1314 5</intersection>
<intersection>1327 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>503.5,1327,507,1327</points>
<connection>
<GID>1420</GID>
<name>IN_4</name></connection>
<intersection>503.5 11</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>478.5,1306.5,491.5,1306.5</points>
<connection>
<GID>1143</GID>
<name>OUT</name></connection>
<intersection>491.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>1757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1295.5,497,1304.5</points>
<intersection>1295.5 1</intersection>
<intersection>1304.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,1295.5,497,1295.5</points>
<connection>
<GID>1144</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1304.5,509,1304.5</points>
<connection>
<GID>1148</GID>
<name>IN_3</name></connection>
<intersection>497 0</intersection>
<intersection>499 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>499,1304.5,499,1313</points>
<intersection>1304.5 2</intersection>
<intersection>1313 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>499,1313,530,1313</points>
<connection>
<GID>1192</GID>
<name>IN_3</name></connection>
<intersection>499 3</intersection>
<intersection>504 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>504,1313,504,1326</points>
<intersection>1313 4</intersection>
<intersection>1326 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>504,1326,507,1326</points>
<connection>
<GID>1420</GID>
<name>IN_3</name></connection>
<intersection>504 5</intersection></hsegment></shape></wire>
<wire>
<ID>1758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1284.5,497,1303.5</points>
<intersection>1284.5 1</intersection>
<intersection>1303.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,1284.5,497,1284.5</points>
<connection>
<GID>1145</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1303.5,509,1303.5</points>
<connection>
<GID>1148</GID>
<name>IN_2</name></connection>
<intersection>497 0</intersection>
<intersection>500 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>500,1303.5,500,1312</points>
<intersection>1303.5 2</intersection>
<intersection>1312 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>500,1312,530,1312</points>
<connection>
<GID>1192</GID>
<name>IN_2</name></connection>
<intersection>500 3</intersection>
<intersection>504.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>504.5,1312,504.5,1325</points>
<intersection>1312 4</intersection>
<intersection>1325 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>504.5,1325,507,1325</points>
<connection>
<GID>1420</GID>
<name>IN_2</name></connection>
<intersection>504.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1274,497,1302.5</points>
<intersection>1274 1</intersection>
<intersection>1302.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>478.5,1274,497,1274</points>
<connection>
<GID>1146</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>497,1302.5,509,1302.5</points>
<connection>
<GID>1148</GID>
<name>IN_1</name></connection>
<intersection>497 0</intersection>
<intersection>501 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>501,1302.5,501,1311</points>
<intersection>1302.5 2</intersection>
<intersection>1311 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>501,1311,530,1311</points>
<connection>
<GID>1192</GID>
<name>IN_1</name></connection>
<intersection>501 3</intersection>
<intersection>505 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>505,1311,505,1324</points>
<intersection>1311 4</intersection>
<intersection>1324 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>505,1324,507,1324</points>
<connection>
<GID>1420</GID>
<name>IN_1</name></connection>
<intersection>505 5</intersection></hsegment></shape></wire>
<wire>
<ID>1760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,1263,497,1301.5</points>
<intersection>1263 2</intersection>
<intersection>1301.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497,1301.5,509,1301.5</points>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection>
<intersection>497 0</intersection>
<intersection>502 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>478.5,1263,497,1263</points>
<connection>
<GID>1147</GID>
<name>OUT</name></connection>
<intersection>497 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>502,1301.5,502,1310</points>
<intersection>1301.5 1</intersection>
<intersection>1310 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>502,1310,530,1310</points>
<connection>
<GID>1192</GID>
<name>IN_0</name></connection>
<intersection>502 3</intersection>
<intersection>505.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>505.5,1310,505.5,1323</points>
<intersection>1310 4</intersection>
<intersection>1323 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>505.5,1323,507,1323</points>
<connection>
<GID>1420</GID>
<name>IN_0</name></connection>
<intersection>505.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1761</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>470,1260,470,1324</points>
<intersection>1260 17</intersection>
<intersection>1324 18</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>470,1260,485,1260</points>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection>
<connection>
<GID>1170</GID>
<name>IN_0</name></connection>
<intersection>470 14</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>454,1324,470,1324</points>
<connection>
<GID>1138</GID>
<name>OUT_0</name></connection>
<intersection>470 14</intersection></hsegment></shape></wire>
<wire>
<ID>1762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,1282,452,1321.5</points>
<intersection>1282 8</intersection>
<intersection>1295 7</intersection>
<intersection>1308.5 6</intersection>
<intersection>1321.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>449,1321.5,452,1321.5</points>
<intersection>449 51</intersection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>449,1308.5,452,1308.5</points>
<intersection>449 50</intersection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>449,1295,452,1295</points>
<intersection>449 49</intersection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>448,1282,452,1282</points>
<intersection>448 53</intersection>
<intersection>449 48</intersection>
<intersection>452 0</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>449,1282,449,1282.5</points>
<connection>
<GID>1103</GID>
<name>clock</name></connection>
<intersection>1282 8</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>449,1295,449,1295.5</points>
<connection>
<GID>1105</GID>
<name>clock</name></connection>
<intersection>1295 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>449,1308.5,449,1309</points>
<connection>
<GID>1136</GID>
<name>clock</name></connection>
<intersection>1308.5 6</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>449,1321.5,449,1322</points>
<connection>
<GID>1138</GID>
<name>clock</name></connection>
<intersection>1321.5 5</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>448,1279,448,1282</points>
<connection>
<GID>1110</GID>
<name>CLK</name></connection>
<intersection>1279 54</intersection>
<intersection>1282 8</intersection></vsegment>
<hsegment>
<ID>54</ID>
<points>448,1279,449,1279</points>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection>
<intersection>448 53</intersection></hsegment></shape></wire>
<wire>
<ID>1763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>476.5,1268,476.5,1346</points>
<connection>
<GID>1147</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1146</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1145</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1144</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1143</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1142</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1141</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1139</GID>
<name>SEL_0</name></connection>
<intersection>1346 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>420.5,1346,476.5,1346</points>
<intersection>420.5 22</intersection>
<intersection>476.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>420.5,1327.5,420.5,1346</points>
<intersection>1327.5 27</intersection>
<intersection>1346 21</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>406,1327.5,420.5,1327.5</points>
<connection>
<GID>1295</GID>
<name>OUT_0</name></connection>
<intersection>408 29</intersection>
<intersection>420.5 22</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>408,1315.5,408,1327.5</points>
<intersection>1315.5 30</intersection>
<intersection>1327.5 27</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>406,1315.5,408,1315.5</points>
<connection>
<GID>1498</GID>
<name>OUT_0</name></connection>
<intersection>408 29</intersection></hsegment></shape></wire>
<wire>
<ID>1764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>475.5,1268,475.5,1345.5</points>
<connection>
<GID>1147</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1146</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1145</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1144</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1143</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1142</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1141</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1139</GID>
<name>SEL_1</name></connection>
<intersection>1345.5 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>420,1345.5,475.5,1345.5</points>
<intersection>420 22</intersection>
<intersection>475.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>420,1328.5,420,1345.5</points>
<intersection>1328.5 25</intersection>
<intersection>1345.5 21</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>408.5,1328.5,420,1328.5</points>
<intersection>408.5 28</intersection>
<intersection>420 22</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>408.5,1316.5,408.5,1328.5</points>
<intersection>1316.5 29</intersection>
<intersection>1328.5 25</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>406,1316.5,408.5,1316.5</points>
<connection>
<GID>1498</GID>
<name>OUT_1</name></connection>
<intersection>408.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>1765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1298.5,491.5,1338</points>
<intersection>1298.5 2</intersection>
<intersection>1338 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1338,491.5,1338</points>
<connection>
<GID>1157</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1298.5,509,1298.5</points>
<connection>
<GID>1172</GID>
<name>IN_7</name></connection>
<intersection>491.5 0</intersection>
<intersection>497.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>497.5,1290,497.5,1298.5</points>
<intersection>1290 4</intersection>
<intersection>1298.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>497.5,1290,530,1290</points>
<connection>
<GID>1194</GID>
<name>IN_7</name></connection>
<intersection>497.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1297.5,491.5,1327</points>
<intersection>1297.5 2</intersection>
<intersection>1327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1327,491.5,1327</points>
<connection>
<GID>1160</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1297.5,509,1297.5</points>
<connection>
<GID>1172</GID>
<name>IN_6</name></connection>
<intersection>491.5 0</intersection>
<intersection>498 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>498,1289,498,1297.5</points>
<intersection>1289 4</intersection>
<intersection>1297.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>498,1289,530,1289</points>
<connection>
<GID>1194</GID>
<name>IN_6</name></connection>
<intersection>498 3</intersection></hsegment></shape></wire>
<wire>
<ID>1767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1296.5,491.5,1316</points>
<intersection>1296.5 2</intersection>
<intersection>1316 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1316,491.5,1316</points>
<connection>
<GID>1162</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1296.5,509,1296.5</points>
<connection>
<GID>1172</GID>
<name>IN_5</name></connection>
<intersection>491.5 0</intersection>
<intersection>500 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>500,1288,500,1296.5</points>
<intersection>1288 4</intersection>
<intersection>1296.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>500,1288,530,1288</points>
<connection>
<GID>1194</GID>
<name>IN_5</name></connection>
<intersection>500 3</intersection></hsegment></shape></wire>
<wire>
<ID>1768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1295.5,491.5,1306.5</points>
<intersection>1295.5 2</intersection>
<intersection>1306.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1306.5,491.5,1306.5</points>
<connection>
<GID>1164</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1295.5,509,1295.5</points>
<connection>
<GID>1172</GID>
<name>IN_4</name></connection>
<intersection>491.5 0</intersection>
<intersection>501.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>501.5,1287,501.5,1295.5</points>
<intersection>1287 4</intersection>
<intersection>1295.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>501.5,1287,530,1287</points>
<connection>
<GID>1194</GID>
<name>IN_4</name></connection>
<intersection>501.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>491.5,1294.5,509,1294.5</points>
<connection>
<GID>1172</GID>
<name>IN_3</name></connection>
<intersection>491.5 2</intersection>
<intersection>503.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>491.5,1294.5,491.5,1295.5</points>
<intersection>1294.5 1</intersection>
<intersection>1295.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>491,1295.5,491.5,1295.5</points>
<connection>
<GID>1165</GID>
<name>OUT</name></connection>
<intersection>491.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>503.5,1286,503.5,1294.5</points>
<intersection>1286 5</intersection>
<intersection>1294.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>503.5,1286,530,1286</points>
<connection>
<GID>1194</GID>
<name>IN_3</name></connection>
<intersection>503.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1770</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1284.5,491.5,1293.5</points>
<intersection>1284.5 1</intersection>
<intersection>1293.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1284.5,491.5,1284.5</points>
<connection>
<GID>1166</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1293.5,509,1293.5</points>
<connection>
<GID>1172</GID>
<name>IN_2</name></connection>
<intersection>491.5 0</intersection>
<intersection>505.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>505.5,1285,505.5,1293.5</points>
<intersection>1285 4</intersection>
<intersection>1293.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>505.5,1285,530,1285</points>
<connection>
<GID>1194</GID>
<name>IN_2</name></connection>
<intersection>505.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1274,491.5,1292.5</points>
<intersection>1274 1</intersection>
<intersection>1292.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491,1274,491.5,1274</points>
<connection>
<GID>1167</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491.5,1292.5,509,1292.5</points>
<connection>
<GID>1172</GID>
<name>IN_1</name></connection>
<intersection>491.5 0</intersection>
<intersection>506.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>506.5,1284,506.5,1292.5</points>
<intersection>1284 4</intersection>
<intersection>1292.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>506.5,1284,530,1284</points>
<connection>
<GID>1194</GID>
<name>IN_1</name></connection>
<intersection>506.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1263,491.5,1291.5</points>
<intersection>1263 2</intersection>
<intersection>1291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>491.5,1291.5,509,1291.5</points>
<connection>
<GID>1172</GID>
<name>IN_0</name></connection>
<intersection>491.5 0</intersection>
<intersection>507.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>491,1263,491.5,1263</points>
<connection>
<GID>1170</GID>
<name>OUT</name></connection>
<intersection>491.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>507.5,1283,507.5,1291.5</points>
<intersection>1283 4</intersection>
<intersection>1291.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>507.5,1283,530,1283</points>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection>
<intersection>507.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,1268,489,1347</points>
<connection>
<GID>1166</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1165</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1164</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1162</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1160</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1157</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1170</GID>
<name>SEL_0</name></connection>
<connection>
<GID>1167</GID>
<name>SEL_0</name></connection>
<intersection>1347 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>421.5,1347,489,1347</points>
<intersection>421.5 25</intersection>
<intersection>489 0</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>421.5,1329.5,421.5,1347</points>
<intersection>1329.5 27</intersection>
<intersection>1347 24</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>409,1329.5,421.5,1329.5</points>
<intersection>409 28</intersection>
<intersection>421.5 25</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>409,1317.5,409,1329.5</points>
<intersection>1317.5 29</intersection>
<intersection>1329.5 27</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>406,1317.5,409,1317.5</points>
<connection>
<GID>1498</GID>
<name>OUT_2</name></connection>
<intersection>409 28</intersection></hsegment></shape></wire>
<wire>
<ID>1774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488,1268,488,1346.5</points>
<connection>
<GID>1166</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1165</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1164</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1162</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1160</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1157</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1170</GID>
<name>SEL_1</name></connection>
<connection>
<GID>1167</GID>
<name>SEL_1</name></connection>
<intersection>1346.5 30</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>421,1346.5,488,1346.5</points>
<intersection>421 31</intersection>
<intersection>488 0</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>421,1330.5,421,1346.5</points>
<intersection>1330.5 33</intersection>
<intersection>1346.5 30</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>409.5,1330.5,421,1330.5</points>
<intersection>409.5 34</intersection>
<intersection>421 31</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>409.5,1318.5,409.5,1330.5</points>
<intersection>1318.5 35</intersection>
<intersection>1330.5 33</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>406,1318.5,409.5,1318.5</points>
<connection>
<GID>1498</GID>
<name>OUT_3</name></connection>
<intersection>409.5 34</intersection></hsegment></shape></wire>
<wire>
<ID>1775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,1291.5,444.5,1331</points>
<intersection>1291.5 1</intersection>
<intersection>1304.5 2</intersection>
<intersection>1318 3</intersection>
<intersection>1331 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,1291.5,446,1291.5</points>
<connection>
<GID>1103</GID>
<name>IN_7</name></connection>
<intersection>444.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444.5,1304.5,446,1304.5</points>
<connection>
<GID>1105</GID>
<name>IN_7</name></connection>
<intersection>444.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>436.5,1318,446,1318</points>
<connection>
<GID>1136</GID>
<name>IN_7</name></connection>
<intersection>436.5 7</intersection>
<intersection>444.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444.5,1331,446,1331</points>
<connection>
<GID>1138</GID>
<name>IN_7</name></connection>
<intersection>444.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>436.5,1281,436.5,1318</points>
<intersection>1281 8</intersection>
<intersection>1318 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>413,1281,436.5,1281</points>
<connection>
<GID>1109</GID>
<name>OUT_7</name></connection>
<intersection>416 9</intersection>
<intersection>436.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>416,1268.5,416,1281</points>
<intersection>1268.5 12</intersection>
<intersection>1281 8</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>415.5,1268.5,416,1268.5</points>
<connection>
<GID>1469</GID>
<name>OUT_7</name></connection>
<intersection>416 9</intersection></hsegment></shape></wire>
<wire>
<ID>1776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,1290.5,444,1330</points>
<intersection>1290.5 4</intersection>
<intersection>1302.5 2</intersection>
<intersection>1303.5 3</intersection>
<intersection>1317 5</intersection>
<intersection>1330 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>437,1302.5,444,1302.5</points>
<intersection>437 7</intersection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>444,1303.5,446,1303.5</points>
<connection>
<GID>1105</GID>
<name>IN_6</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>444,1290.5,446,1290.5</points>
<connection>
<GID>1103</GID>
<name>IN_6</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>444,1317,446,1317</points>
<connection>
<GID>1136</GID>
<name>IN_6</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>444,1330,446,1330</points>
<connection>
<GID>1138</GID>
<name>IN_6</name></connection>
<intersection>444 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>437,1280,437,1302.5</points>
<intersection>1280 8</intersection>
<intersection>1302.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>413,1280,437,1280</points>
<connection>
<GID>1109</GID>
<name>OUT_6</name></connection>
<intersection>416.5 9</intersection>
<intersection>437 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>416.5,1267.5,416.5,1280</points>
<intersection>1267.5 10</intersection>
<intersection>1280 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>415.5,1267.5,416.5,1267.5</points>
<connection>
<GID>1469</GID>
<name>OUT_6</name></connection>
<intersection>416.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>1777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443.5,1289.5,443.5,1329</points>
<intersection>1289.5 5</intersection>
<intersection>1300.5 2</intersection>
<intersection>1302.5 4</intersection>
<intersection>1316 3</intersection>
<intersection>1329 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>437.5,1300.5,443.5,1300.5</points>
<intersection>437.5 7</intersection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>443.5,1316,446,1316</points>
<connection>
<GID>1136</GID>
<name>IN_5</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>443.5,1302.5,446,1302.5</points>
<connection>
<GID>1105</GID>
<name>IN_5</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>443.5,1289.5,446,1289.5</points>
<connection>
<GID>1103</GID>
<name>IN_5</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443.5,1329,446,1329</points>
<connection>
<GID>1138</GID>
<name>IN_5</name></connection>
<intersection>443.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>437.5,1279,437.5,1300.5</points>
<intersection>1279 8</intersection>
<intersection>1300.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>413,1279,437.5,1279</points>
<connection>
<GID>1109</GID>
<name>OUT_5</name></connection>
<intersection>417 9</intersection>
<intersection>437.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>417,1266.5,417,1279</points>
<intersection>1266.5 10</intersection>
<intersection>1279 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>415.5,1266.5,417,1266.5</points>
<connection>
<GID>1469</GID>
<name>OUT_5</name></connection>
<intersection>417 9</intersection></hsegment></shape></wire>
<wire>
<ID>1778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443,1288.5,443,1328</points>
<intersection>1288.5 5</intersection>
<intersection>1298.5 2</intersection>
<intersection>1301.5 4</intersection>
<intersection>1315 3</intersection>
<intersection>1328 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>438,1298.5,443,1298.5</points>
<intersection>438 7</intersection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>443,1315,446,1315</points>
<connection>
<GID>1136</GID>
<name>IN_4</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>443,1301.5,446,1301.5</points>
<connection>
<GID>1105</GID>
<name>IN_4</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>443,1288.5,446,1288.5</points>
<connection>
<GID>1103</GID>
<name>IN_4</name></connection>
<intersection>443 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>443,1328,446,1328</points>
<connection>
<GID>1138</GID>
<name>IN_4</name></connection>
<intersection>443 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>438,1278,438,1298.5</points>
<intersection>1278 8</intersection>
<intersection>1298.5 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>413,1278,438,1278</points>
<connection>
<GID>1109</GID>
<name>OUT_4</name></connection>
<intersection>417.5 9</intersection>
<intersection>438 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>417.5,1265.5,417.5,1278</points>
<intersection>1265.5 10</intersection>
<intersection>1278 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>415.5,1265.5,417.5,1265.5</points>
<connection>
<GID>1469</GID>
<name>OUT_4</name></connection>
<intersection>417.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>1779</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442.5,1287.5,442.5,1327</points>
<intersection>1287.5 4</intersection>
<intersection>1291 2</intersection>
<intersection>1300.5 3</intersection>
<intersection>1314 12</intersection>
<intersection>1327 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>438.5,1291,442.5,1291</points>
<intersection>438.5 10</intersection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>442.5,1300.5,446,1300.5</points>
<connection>
<GID>1105</GID>
<name>IN_3</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>442.5,1287.5,446,1287.5</points>
<connection>
<GID>1103</GID>
<name>IN_3</name></connection>
<intersection>442.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>442.5,1327,446,1327</points>
<connection>
<GID>1138</GID>
<name>IN_3</name></connection>
<intersection>442.5 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>438.5,1277,438.5,1291</points>
<intersection>1277 11</intersection>
<intersection>1291 2</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>413,1277,438.5,1277</points>
<connection>
<GID>1109</GID>
<name>OUT_3</name></connection>
<intersection>418 13</intersection>
<intersection>438.5 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>442.5,1314,446,1314</points>
<connection>
<GID>1136</GID>
<name>IN_3</name></connection>
<intersection>442.5 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>418,1264.5,418,1277</points>
<intersection>1264.5 14</intersection>
<intersection>1277 11</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>415.5,1264.5,418,1264.5</points>
<connection>
<GID>1469</GID>
<name>OUT_3</name></connection>
<intersection>418 13</intersection></hsegment></shape></wire>
<wire>
<ID>1780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442,1286.5,442,1326</points>
<intersection>1286.5 1</intersection>
<intersection>1289 2</intersection>
<intersection>1299.5 3</intersection>
<intersection>1313 4</intersection>
<intersection>1326 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,1286.5,446,1286.5</points>
<connection>
<GID>1103</GID>
<name>IN_2</name></connection>
<intersection>442 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>439,1289,442,1289</points>
<intersection>439 6</intersection>
<intersection>442 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>442,1299.5,446,1299.5</points>
<connection>
<GID>1105</GID>
<name>IN_2</name></connection>
<intersection>442 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>442,1313,446,1313</points>
<connection>
<GID>1136</GID>
<name>IN_2</name></connection>
<intersection>442 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>442,1326,446,1326</points>
<connection>
<GID>1138</GID>
<name>IN_2</name></connection>
<intersection>442 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>439,1276,439,1289</points>
<intersection>1276 7</intersection>
<intersection>1289 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>413,1276,439,1276</points>
<connection>
<GID>1109</GID>
<name>OUT_2</name></connection>
<intersection>418.5 8</intersection>
<intersection>439 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>418.5,1263.5,418.5,1276</points>
<intersection>1263.5 9</intersection>
<intersection>1276 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>415.5,1263.5,418.5,1263.5</points>
<connection>
<GID>1469</GID>
<name>OUT_2</name></connection>
<intersection>418.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,1285.5,441.5,1325</points>
<intersection>1285.5 1</intersection>
<intersection>1287 2</intersection>
<intersection>1298.5 3</intersection>
<intersection>1312 4</intersection>
<intersection>1325 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>441.5,1285.5,446,1285.5</points>
<connection>
<GID>1103</GID>
<name>IN_1</name></connection>
<intersection>441.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>439.5,1287,441.5,1287</points>
<intersection>439.5 6</intersection>
<intersection>441.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>441.5,1298.5,446,1298.5</points>
<connection>
<GID>1105</GID>
<name>IN_1</name></connection>
<intersection>441.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>441.5,1312,446,1312</points>
<connection>
<GID>1136</GID>
<name>IN_1</name></connection>
<intersection>441.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>441.5,1325,446,1325</points>
<connection>
<GID>1138</GID>
<name>IN_1</name></connection>
<intersection>441.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>439.5,1275,439.5,1287</points>
<intersection>1275 7</intersection>
<intersection>1287 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>413,1275,439.5,1275</points>
<connection>
<GID>1109</GID>
<name>OUT_1</name></connection>
<intersection>419 8</intersection>
<intersection>439.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>419,1262.5,419,1275</points>
<intersection>1262.5 9</intersection>
<intersection>1275 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>415.5,1262.5,419,1262.5</points>
<connection>
<GID>1469</GID>
<name>OUT_1</name></connection>
<intersection>419 8</intersection></hsegment></shape></wire>
<wire>
<ID>1782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441,1285,441,1324</points>
<intersection>1285 1</intersection>
<intersection>1297.5 3</intersection>
<intersection>1311 4</intersection>
<intersection>1324 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>440,1285,446,1285</points>
<intersection>440 6</intersection>
<intersection>441 0</intersection>
<intersection>446 11</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>441,1297.5,446,1297.5</points>
<connection>
<GID>1105</GID>
<name>IN_0</name></connection>
<intersection>441 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>441,1311,446,1311</points>
<connection>
<GID>1136</GID>
<name>IN_0</name></connection>
<intersection>441 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>441,1324,446,1324</points>
<connection>
<GID>1138</GID>
<name>IN_0</name></connection>
<intersection>441 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>440,1274,440,1285</points>
<intersection>1274 7</intersection>
<intersection>1285 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>413,1274,440,1274</points>
<connection>
<GID>1109</GID>
<name>OUT_0</name></connection>
<intersection>419.5 12</intersection>
<intersection>440 6</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>446,1284.5,446,1285</points>
<connection>
<GID>1103</GID>
<name>IN_0</name></connection>
<intersection>1285 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>419.5,1261.5,419.5,1274</points>
<intersection>1261.5 13</intersection>
<intersection>1274 7</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>415.5,1261.5,419.5,1261.5</points>
<connection>
<GID>1469</GID>
<name>OUT_0</name></connection>
<intersection>419.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>1783</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>706.5,1335,707,1335</points>
<connection>
<GID>1333</GID>
<name>IN_0</name></connection>
<intersection>706.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>706.5,1334.5,706.5,1335</points>
<connection>
<GID>1179</GID>
<name>OUT_1</name></connection>
<intersection>1335 1</intersection></vsegment></shape></wire>
<wire>
<ID>1784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532,1291.5,532,1292.5</points>
<connection>
<GID>1194</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1205</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1785</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>454.5,1341,485,1341</points>
<connection>
<GID>1157</GID>
<name>IN_3</name></connection>
<connection>
<GID>1139</GID>
<name>IN_3</name></connection>
<intersection>454.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>454.5,1291.5,454.5,1341</points>
<intersection>1291.5 5</intersection>
<intersection>1341 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1291.5,454.5,1291.5</points>
<connection>
<GID>1103</GID>
<name>OUT_7</name></connection>
<intersection>454.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>591.5,1353.5,591.5,1386.5</points>
<connection>
<GID>1125</GID>
<name>ENABLE_0</name></connection>
<intersection>1379.5 2</intersection>
<intersection>1386.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,1386.5,591.5,1386.5</points>
<connection>
<GID>1107</GID>
<name>ENABLE_0</name></connection>
<intersection>591.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>591.5,1379.5,597,1379.5</points>
<connection>
<GID>1286</GID>
<name>OUT_0</name></connection>
<intersection>591.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1788</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1311,570.5,1311</points>
<connection>
<GID>1289</GID>
<name>IN_5</name></connection>
<intersection>536 7</intersection>
<intersection>566 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>566,1288,566,1311</points>
<intersection>1288 4</intersection>
<intersection>1311 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>566,1288,570.5,1288</points>
<connection>
<GID>1290</GID>
<name>IN_5</name></connection>
<intersection>566 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>536,1311,536,1312</points>
<intersection>1311 1</intersection>
<intersection>1312 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>534,1312,536,1312</points>
<connection>
<GID>1192</GID>
<name>OUT_2</name></connection>
<intersection>536 7</intersection></hsegment></shape></wire>
<wire>
<ID>1789</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>535.5,1309,570.5,1309</points>
<connection>
<GID>1289</GID>
<name>IN_3</name></connection>
<intersection>535.5 5</intersection>
<intersection>567 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>567,1286,567,1309</points>
<intersection>1286 4</intersection>
<intersection>1309 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>567,1286,570.5,1286</points>
<connection>
<GID>1290</GID>
<name>IN_3</name></connection>
<intersection>567 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>535.5,1309,535.5,1311</points>
<intersection>1309 1</intersection>
<intersection>1311 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1311,535.5,1311</points>
<connection>
<GID>1192</GID>
<name>OUT_1</name></connection>
<intersection>535.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1790</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>535,1307,570.5,1307</points>
<connection>
<GID>1289</GID>
<name>IN_1</name></connection>
<intersection>535 5</intersection>
<intersection>568 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>568,1284,568,1307</points>
<intersection>1284 4</intersection>
<intersection>1307 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>568,1284,570.5,1284</points>
<connection>
<GID>1290</GID>
<name>IN_1</name></connection>
<intersection>568 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>535,1307,535,1310</points>
<intersection>1307 1</intersection>
<intersection>1310 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1310,535,1310</points>
<connection>
<GID>1192</GID>
<name>OUT_0</name></connection>
<intersection>535 5</intersection></hsegment></shape></wire>
<wire>
<ID>1791</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534,1297,570.5,1297</points>
<connection>
<GID>1290</GID>
<name>IN_14</name></connection>
<intersection>534 5</intersection>
<intersection>561.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>561.5,1297,561.5,1320</points>
<intersection>1297 1</intersection>
<intersection>1320 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>561.5,1320,570.5,1320</points>
<connection>
<GID>1289</GID>
<name>IN_14</name></connection>
<intersection>561.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>534,1290,534,1297</points>
<connection>
<GID>1194</GID>
<name>OUT_7</name></connection>
<intersection>1297 1</intersection></vsegment></shape></wire>
<wire>
<ID>1792</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534.5,1295,570.5,1295</points>
<connection>
<GID>1290</GID>
<name>IN_12</name></connection>
<intersection>534.5 5</intersection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>562.5,1295,562.5,1318</points>
<intersection>1295 1</intersection>
<intersection>1318 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>562.5,1318,570.5,1318</points>
<connection>
<GID>1289</GID>
<name>IN_12</name></connection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>534.5,1289,534.5,1295</points>
<intersection>1289 6</intersection>
<intersection>1295 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1289,534.5,1289</points>
<connection>
<GID>1194</GID>
<name>OUT_6</name></connection>
<intersection>534.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1793</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>535,1293,570.5,1293</points>
<connection>
<GID>1290</GID>
<name>IN_10</name></connection>
<intersection>535 5</intersection>
<intersection>563.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>563.5,1293,563.5,1316</points>
<intersection>1293 1</intersection>
<intersection>1316 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>563.5,1316,570.5,1316</points>
<connection>
<GID>1289</GID>
<name>IN_10</name></connection>
<intersection>563.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>535,1288,535,1293</points>
<intersection>1288 6</intersection>
<intersection>1293 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1288,535,1288</points>
<connection>
<GID>1194</GID>
<name>OUT_5</name></connection>
<intersection>535 5</intersection></hsegment></shape></wire>
<wire>
<ID>1794</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>535.5,1291,570.5,1291</points>
<connection>
<GID>1290</GID>
<name>IN_8</name></connection>
<intersection>535.5 5</intersection>
<intersection>564.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>564.5,1291,564.5,1314</points>
<intersection>1291 1</intersection>
<intersection>1314 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>564.5,1314,570.5,1314</points>
<connection>
<GID>1289</GID>
<name>IN_8</name></connection>
<intersection>564.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>535.5,1287,535.5,1291</points>
<intersection>1287 6</intersection>
<intersection>1291 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1287,535.5,1287</points>
<connection>
<GID>1194</GID>
<name>OUT_4</name></connection>
<intersection>535.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1795</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536,1289,570.5,1289</points>
<connection>
<GID>1290</GID>
<name>IN_6</name></connection>
<intersection>536 5</intersection>
<intersection>565.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>565.5,1289,565.5,1312</points>
<intersection>1289 1</intersection>
<intersection>1312 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>565.5,1312,570.5,1312</points>
<connection>
<GID>1289</GID>
<name>IN_6</name></connection>
<intersection>565.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>536,1286,536,1289</points>
<intersection>1286 6</intersection>
<intersection>1289 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1286,536,1286</points>
<connection>
<GID>1194</GID>
<name>OUT_3</name></connection>
<intersection>536 5</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>671,1361,671.5,1361</points>
<connection>
<GID>847</GID>
<name>OUT</name></connection>
<connection>
<GID>969</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1796</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>536.5,1287,570.5,1287</points>
<connection>
<GID>1290</GID>
<name>IN_4</name></connection>
<intersection>536.5 5</intersection>
<intersection>566.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>566.5,1287,566.5,1310</points>
<intersection>1287 1</intersection>
<intersection>1310 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>566.5,1310,570.5,1310</points>
<connection>
<GID>1289</GID>
<name>IN_4</name></connection>
<intersection>566.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>536.5,1285,536.5,1287</points>
<intersection>1285 6</intersection>
<intersection>1287 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1285,536.5,1285</points>
<connection>
<GID>1194</GID>
<name>OUT_2</name></connection>
<intersection>536.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>710.5,1296,710.5,1297.5</points>
<connection>
<GID>841</GID>
<name>OUT_0</name></connection>
<intersection>1296 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>710.5,1296,711.5,1296</points>
<connection>
<GID>1075</GID>
<name>ENABLE</name></connection>
<intersection>710.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1797</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>537,1285,570.5,1285</points>
<connection>
<GID>1290</GID>
<name>IN_2</name></connection>
<intersection>537 5</intersection>
<intersection>567.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>567.5,1285,567.5,1308</points>
<intersection>1285 1</intersection>
<intersection>1308 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>567.5,1308,570.5,1308</points>
<connection>
<GID>1289</GID>
<name>IN_2</name></connection>
<intersection>567.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>537,1284,537,1285</points>
<intersection>1284 6</intersection>
<intersection>1285 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>534,1284,537,1284</points>
<connection>
<GID>1194</GID>
<name>OUT_1</name></connection>
<intersection>537 5</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>659,1344,659,1344</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<connection>
<GID>1296</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1798</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534,1283,570.5,1283</points>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection>
<connection>
<GID>1194</GID>
<name>OUT_0</name></connection>
<intersection>568.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>568.5,1283,568.5,1306</points>
<intersection>1283 1</intersection>
<intersection>1306 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>568.5,1306,570.5,1306</points>
<connection>
<GID>1289</GID>
<name>IN_0</name></connection>
<intersection>568.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>659,1338.5,659,1338.5</points>
<connection>
<GID>976</GID>
<name>IN_0</name></connection>
<connection>
<GID>1052</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1799</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1283,585.5,1283</points>
<connection>
<GID>1134</GID>
<name>IN_0</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1307.5,680.5,1311.5</points>
<connection>
<GID>968</GID>
<name>IN_0</name></connection>
<intersection>1307.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1307.5,692,1307.5</points>
<connection>
<GID>990</GID>
<name>IN_7</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1800</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1285,585.5,1285</points>
<connection>
<GID>1134</GID>
<name>IN_2</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1801</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1284,585.5,1284</points>
<connection>
<GID>1134</GID>
<name>IN_1</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1802</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1286,585.5,1286</points>
<connection>
<GID>1134</GID>
<name>IN_3</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1309.5,680.5,1313.5</points>
<connection>
<GID>970</GID>
<name>IN_0</name></connection>
<intersection>1309.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1309.5,692,1309.5</points>
<connection>
<GID>990</GID>
<name>IN_9</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1803</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1287,585.5,1287</points>
<connection>
<GID>1134</GID>
<name>IN_4</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1311.5,680.5,1315.5</points>
<connection>
<GID>971</GID>
<name>IN_0</name></connection>
<intersection>1311.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1311.5,692,1311.5</points>
<connection>
<GID>990</GID>
<name>IN_11</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1804</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1288,585.5,1288</points>
<connection>
<GID>1134</GID>
<name>IN_5</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1805</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1290,585.5,1290</points>
<connection>
<GID>1134</GID>
<name>IN_7</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1806</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1289,585.5,1289</points>
<connection>
<GID>1134</GID>
<name>IN_6</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1807</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1292,585.5,1292</points>
<connection>
<GID>1134</GID>
<name>IN_9</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1808</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1293,585.5,1293</points>
<connection>
<GID>1134</GID>
<name>IN_10</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1809</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1291,585.5,1291</points>
<connection>
<GID>1134</GID>
<name>IN_8</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1810</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1294,585.5,1294</points>
<connection>
<GID>1134</GID>
<name>IN_11</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1303.5,680.5,1307.5</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<intersection>1303.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1303.5,692,1303.5</points>
<connection>
<GID>990</GID>
<name>IN_3</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1811</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1295,585.5,1295</points>
<connection>
<GID>1134</GID>
<name>IN_12</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1812</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1297,585.5,1297</points>
<connection>
<GID>1134</GID>
<name>IN_14</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,1344,432,1344</points>
<connection>
<GID>1181</GID>
<name>ENABLE</name></connection>
<connection>
<GID>1002</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1813</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1296,585.5,1296</points>
<connection>
<GID>1134</GID>
<name>IN_13</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1814</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1298,585.5,1298</points>
<connection>
<GID>1134</GID>
<name>IN_15</name></connection>
<connection>
<GID>1290</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1815</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1307,585.5,1307</points>
<connection>
<GID>1133</GID>
<name>IN_1</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1816</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1310,585.5,1310</points>
<connection>
<GID>1133</GID>
<name>IN_4</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1817</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1311,585.5,1311</points>
<connection>
<GID>1133</GID>
<name>IN_5</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1818</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1309,585.5,1309</points>
<connection>
<GID>1133</GID>
<name>IN_3</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1819</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1308,585.5,1308</points>
<connection>
<GID>1133</GID>
<name>IN_2</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1820</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1312,585.5,1312</points>
<connection>
<GID>1133</GID>
<name>IN_6</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1821</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1313,585.5,1313</points>
<connection>
<GID>1133</GID>
<name>IN_7</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1822</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1306,585.5,1306</points>
<connection>
<GID>1133</GID>
<name>IN_0</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1823</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1319,585.5,1319</points>
<connection>
<GID>1133</GID>
<name>IN_13</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1824</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1315,585.5,1315</points>
<connection>
<GID>1133</GID>
<name>IN_9</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1315.5,680.5,1319.5</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<intersection>1315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1315.5,692,1315.5</points>
<connection>
<GID>990</GID>
<name>IN_15</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1825</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1318,585.5,1318</points>
<connection>
<GID>1133</GID>
<name>IN_12</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1057</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,1338,533,1345</points>
<intersection>1338 1</intersection>
<intersection>1345 12</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>529,1338,533,1338</points>
<connection>
<GID>1005</GID>
<name>IN_0</name></connection>
<intersection>533 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>533,1345,558,1345</points>
<connection>
<GID>1015</GID>
<name>IN_0</name></connection>
<intersection>533 0</intersection></hsegment></shape></wire>
<wire>
<ID>1826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1320,585.5,1320</points>
<connection>
<GID>1133</GID>
<name>IN_14</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1827</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1316,585.5,1316</points>
<connection>
<GID>1133</GID>
<name>IN_10</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1828</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1317,585.5,1317</points>
<connection>
<GID>1133</GID>
<name>IN_11</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1314,585.5,1314</points>
<connection>
<GID>1133</GID>
<name>IN_8</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>529,1352,558,1352</points>
<connection>
<GID>1015</GID>
<name>IN_7</name></connection>
<connection>
<GID>1014</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1830</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>574.5,1321,585.5,1321</points>
<connection>
<GID>1133</GID>
<name>IN_15</name></connection>
<connection>
<GID>1289</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1831</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>553.5,1390.5,553.5,1405.5</points>
<intersection>1390.5 3</intersection>
<intersection>1405.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>553.5,1405.5,557,1405.5</points>
<connection>
<GID>1220</GID>
<name>IN_0</name></connection>
<intersection>553.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>553,1390.5,553.5,1390.5</points>
<connection>
<GID>1102</GID>
<name>OUT_7</name></connection>
<intersection>553.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1832</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>554,1389.5,554,1403.5</points>
<intersection>1389.5 3</intersection>
<intersection>1403.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>554,1403.5,557,1403.5</points>
<connection>
<GID>1221</GID>
<name>IN_0</name></connection>
<intersection>554 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>553,1389.5,554,1389.5</points>
<connection>
<GID>1102</GID>
<name>OUT_6</name></connection>
<intersection>554 1</intersection></hsegment></shape></wire>
<wire>
<ID>1833</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>554.5,1388.5,554.5,1401.5</points>
<intersection>1388.5 3</intersection>
<intersection>1401.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>554.5,1401.5,557,1401.5</points>
<connection>
<GID>1223</GID>
<name>IN_0</name></connection>
<intersection>554.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>553,1388.5,554.5,1388.5</points>
<connection>
<GID>1102</GID>
<name>OUT_5</name></connection>
<intersection>554.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1834</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>555,1387.5,555,1399.5</points>
<intersection>1387.5 4</intersection>
<intersection>1399.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>553,1387.5,555,1387.5</points>
<connection>
<GID>1102</GID>
<name>OUT_4</name></connection>
<intersection>555 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>555,1399.5,557,1399.5</points>
<connection>
<GID>1226</GID>
<name>IN_0</name></connection>
<intersection>555 1</intersection></hsegment></shape></wire>
<wire>
<ID>1835</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>555.5,1386.5,555.5,1397.5</points>
<intersection>1386.5 4</intersection>
<intersection>1397.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>553,1386.5,555.5,1386.5</points>
<connection>
<GID>1102</GID>
<name>OUT_3</name></connection>
<intersection>555.5 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>555.5,1397.5,557,1397.5</points>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection>
<intersection>555.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1836</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>556,1385.5,556,1395.5</points>
<intersection>1385.5 4</intersection>
<intersection>1395.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>553,1385.5,556,1385.5</points>
<connection>
<GID>1102</GID>
<name>OUT_2</name></connection>
<intersection>556 1</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>556,1395.5,557,1395.5</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<intersection>556 1</intersection></hsegment></shape></wire>
<wire>
<ID>1837</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>706.5,1333,707,1333</points>
<connection>
<GID>1357</GID>
<name>IN_0</name></connection>
<intersection>706.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>706.5,1333,706.5,1333.5</points>
<connection>
<GID>1179</GID>
<name>OUT_2</name></connection>
<intersection>1333 3</intersection></vsegment></shape></wire>
<wire>
<ID>1838</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>557,1383.5,557,1391.5</points>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection>
<intersection>1383.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>553,1383.5,557,1383.5</points>
<connection>
<GID>1102</GID>
<name>OUT_0</name></connection>
<intersection>557 1</intersection></hsegment></shape></wire>
<wire>
<ID>1839</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>421,1365.5,428,1365.5</points>
<connection>
<GID>1235</GID>
<name>IN_7</name></connection>
<connection>
<GID>1236</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1840</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>421.5,1364.5,428,1364.5</points>
<connection>
<GID>1235</GID>
<name>IN_6</name></connection>
<intersection>421.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>421.5,1363.5,421.5,1364.5</points>
<intersection>1363.5 4</intersection>
<intersection>1364.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>421,1363.5,421.5,1363.5</points>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection>
<intersection>421.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1841</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>421,1359.5,422.5,1359.5</points>
<connection>
<GID>1239</GID>
<name>IN_0</name></connection>
<intersection>422.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>422.5,1359.5,422.5,1362.5</points>
<intersection>1359.5 1</intersection>
<intersection>1362.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>422.5,1362.5,428,1362.5</points>
<connection>
<GID>1235</GID>
<name>IN_4</name></connection>
<intersection>422.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1844</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424,1353.5,424,1359.5</points>
<intersection>1353.5 5</intersection>
<intersection>1359.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>421,1353.5,424,1353.5</points>
<connection>
<GID>1242</GID>
<name>IN_0</name></connection>
<intersection>424 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>424,1359.5,428,1359.5</points>
<connection>
<GID>1235</GID>
<name>IN_1</name></connection>
<intersection>424 0</intersection></hsegment></shape></wire>
<wire>
<ID>1845</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,1351.5,424.5,1358.5</points>
<intersection>1351.5 5</intersection>
<intersection>1358.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>424.5,1358.5,428,1358.5</points>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>421,1351.5,424.5,1351.5</points>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1846</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509,1331.5,509,1332.5</points>
<connection>
<GID>1420</GID>
<name>ENABLE_0</name></connection>
<intersection>1332.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>507.5,1332.5,509,1332.5</points>
<connection>
<GID>1435</GID>
<name>IN_0</name></connection>
<intersection>509 0</intersection></hsegment></shape></wire>
<wire>
<ID>1847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>542,1323,542,1335</points>
<intersection>1323 1</intersection>
<intersection>1335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1323,542,1323</points>
<connection>
<GID>1420</GID>
<name>OUT_0</name></connection>
<intersection>542 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>542,1335,589.5,1335</points>
<connection>
<GID>1439</GID>
<name>IN_0</name></connection>
<intersection>542 0</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>530,1351,558,1351</points>
<connection>
<GID>1015</GID>
<name>IN_6</name></connection>
<intersection>530 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>530,1350,530,1351</points>
<intersection>1350 13</intersection>
<intersection>1351 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>529,1350,530,1350</points>
<connection>
<GID>1013</GID>
<name>IN_0</name></connection>
<intersection>530 8</intersection></hsegment></shape></wire>
<wire>
<ID>1848</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1366,445,1366</points>
<connection>
<GID>1244</GID>
<name>IN_7</name></connection>
<intersection>432 15</intersection>
<intersection>441.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>441.5,1366,441.5,1381</points>
<intersection>1366 1</intersection>
<intersection>1381 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>432,1381,441.5,1381</points>
<connection>
<GID>1302</GID>
<name>OUT_7</name></connection>
<intersection>441.5 6</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>432,1365.5,432,1366</points>
<connection>
<GID>1235</GID>
<name>OUT_7</name></connection>
<intersection>1366 1</intersection></vsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>530.5,1350,558,1350</points>
<connection>
<GID>1015</GID>
<name>IN_5</name></connection>
<intersection>530.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>530.5,1348,530.5,1350</points>
<intersection>1348 16</intersection>
<intersection>1350 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>529,1348,530.5,1348</points>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection>
<intersection>530.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>1849</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432,1365,445,1365</points>
<connection>
<GID>1244</GID>
<name>IN_6</name></connection>
<intersection>432 13</intersection>
<intersection>441 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>441,1365,441,1380</points>
<intersection>1365 2</intersection>
<intersection>1380 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1380,441,1380</points>
<connection>
<GID>1302</GID>
<name>OUT_6</name></connection>
<intersection>441 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1364.5,432,1365</points>
<connection>
<GID>1235</GID>
<name>OUT_6</name></connection>
<intersection>1365 2</intersection></vsegment></shape></wire>
<wire>
<ID>1850</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1364,445,1364</points>
<connection>
<GID>1244</GID>
<name>IN_5</name></connection>
<intersection>432 13</intersection>
<intersection>440.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>440.5,1364,440.5,1379</points>
<intersection>1364 1</intersection>
<intersection>1379 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1379,440.5,1379</points>
<connection>
<GID>1302</GID>
<name>OUT_5</name></connection>
<intersection>440.5 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1363.5,432,1364</points>
<connection>
<GID>1235</GID>
<name>OUT_5</name></connection>
<intersection>1364 1</intersection></vsegment></shape></wire>
<wire>
<ID>1851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1363,445,1363</points>
<connection>
<GID>1244</GID>
<name>IN_4</name></connection>
<intersection>432 13</intersection>
<intersection>440 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>440,1363,440,1378</points>
<intersection>1363 1</intersection>
<intersection>1378 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1378,440,1378</points>
<connection>
<GID>1302</GID>
<name>OUT_4</name></connection>
<intersection>440 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1362.5,432,1363</points>
<connection>
<GID>1235</GID>
<name>OUT_4</name></connection>
<intersection>1363 1</intersection></vsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>531,1349,558,1349</points>
<connection>
<GID>1015</GID>
<name>IN_4</name></connection>
<intersection>531 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>531,1346,531,1349</points>
<intersection>1346 7</intersection>
<intersection>1349 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>529,1346,531,1346</points>
<connection>
<GID>1009</GID>
<name>IN_0</name></connection>
<intersection>531 3</intersection></hsegment></shape></wire>
<wire>
<ID>1852</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1362,445,1362</points>
<connection>
<GID>1244</GID>
<name>IN_3</name></connection>
<intersection>432 13</intersection>
<intersection>439.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>439.5,1362,439.5,1377</points>
<intersection>1362 1</intersection>
<intersection>1377 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1377,439.5,1377</points>
<connection>
<GID>1302</GID>
<name>OUT_3</name></connection>
<intersection>439.5 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1361.5,432,1362</points>
<connection>
<GID>1235</GID>
<name>OUT_3</name></connection>
<intersection>1362 1</intersection></vsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531.5,1344,531.5,1348</points>
<intersection>1344 2</intersection>
<intersection>1348 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>531.5,1348,558,1348</points>
<connection>
<GID>1015</GID>
<name>IN_3</name></connection>
<intersection>531.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,1344,531.5,1344</points>
<connection>
<GID>1008</GID>
<name>IN_0</name></connection>
<intersection>531.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1853</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>432,1361,445,1361</points>
<connection>
<GID>1244</GID>
<name>IN_2</name></connection>
<intersection>432 13</intersection>
<intersection>439 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>439,1361,439,1376</points>
<intersection>1361 2</intersection>
<intersection>1376 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1376,439,1376</points>
<connection>
<GID>1302</GID>
<name>OUT_2</name></connection>
<intersection>439 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1360.5,432,1361</points>
<connection>
<GID>1235</GID>
<name>OUT_2</name></connection>
<intersection>1361 2</intersection></vsegment></shape></wire>
<wire>
<ID>1854</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1360,445,1360</points>
<connection>
<GID>1244</GID>
<name>IN_1</name></connection>
<intersection>432 13</intersection>
<intersection>438.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>438.5,1360,438.5,1375</points>
<intersection>1360 1</intersection>
<intersection>1375 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>432,1375,438.5,1375</points>
<connection>
<GID>1302</GID>
<name>OUT_1</name></connection>
<intersection>438.5 4</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>432,1359.5,432,1360</points>
<connection>
<GID>1235</GID>
<name>OUT_1</name></connection>
<intersection>1360 1</intersection></vsegment></shape></wire>
<wire>
<ID>1855</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,1359,445,1359</points>
<connection>
<GID>1244</GID>
<name>IN_0</name></connection>
<intersection>432 15</intersection>
<intersection>438 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>438,1359,438,1374</points>
<intersection>1359 1</intersection>
<intersection>1374 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>432,1374,438,1374</points>
<connection>
<GID>1302</GID>
<name>OUT_0</name></connection>
<intersection>438 4</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>432,1358.5,432,1359</points>
<connection>
<GID>1235</GID>
<name>OUT_0</name></connection>
<intersection>1359 1</intersection></vsegment></shape></wire>
<wire>
<ID>1856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422,1361.5,422,1363.5</points>
<intersection>1361.5 3</intersection>
<intersection>1363.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>422,1363.5,428,1363.5</points>
<connection>
<GID>1235</GID>
<name>IN_5</name></connection>
<intersection>422 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>421,1361.5,422,1361.5</points>
<connection>
<GID>1238</GID>
<name>IN_0</name></connection>
<intersection>422 0</intersection></hsegment></shape></wire>
<wire>
<ID>1857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538.5,1330,538.5,1342</points>
<intersection>1330 1</intersection>
<intersection>1342 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1330,538.5,1330</points>
<connection>
<GID>1420</GID>
<name>OUT_7</name></connection>
<intersection>538.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538.5,1342,589.5,1342</points>
<connection>
<GID>1439</GID>
<name>IN_7</name></connection>
<intersection>538.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1858</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>451.5,1373,455,1373</points>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection>
<intersection>451.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>451.5,1366,451.5,1373</points>
<intersection>1366 16</intersection>
<intersection>1373 3</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>449,1366,451.5,1366</points>
<connection>
<GID>1244</GID>
<name>OUT_7</name></connection>
<intersection>451.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>1859</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,1365,452,1371</points>
<intersection>1365 3</intersection>
<intersection>1371 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452,1371,455,1371</points>
<connection>
<GID>1249</GID>
<name>IN_0</name></connection>
<intersection>452 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>449,1365,452,1365</points>
<connection>
<GID>1244</GID>
<name>OUT_6</name></connection>
<intersection>452 0</intersection></hsegment></shape></wire>
<wire>
<ID>1860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,1364,452.5,1369</points>
<intersection>1364 3</intersection>
<intersection>1369 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,1369,455,1369</points>
<connection>
<GID>1250</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>449,1364,452.5,1364</points>
<connection>
<GID>1244</GID>
<name>OUT_5</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1861</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453,1363,453,1367</points>
<intersection>1363 3</intersection>
<intersection>1367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453,1367,455,1367</points>
<connection>
<GID>1251</GID>
<name>IN_0</name></connection>
<intersection>453 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>449,1363,453,1363</points>
<connection>
<GID>1244</GID>
<name>OUT_4</name></connection>
<intersection>453 0</intersection></hsegment></shape></wire>
<wire>
<ID>1862</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>453.5,1362,453.5,1365</points>
<intersection>1362 3</intersection>
<intersection>1365 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>453.5,1365,455,1365</points>
<connection>
<GID>1252</GID>
<name>IN_0</name></connection>
<intersection>453.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>449,1362,453.5,1362</points>
<connection>
<GID>1244</GID>
<name>OUT_3</name></connection>
<intersection>453.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1863</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,1361,454,1361</points>
<connection>
<GID>1244</GID>
<name>OUT_2</name></connection>
<intersection>454 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>454,1361,454,1363</points>
<intersection>1361 1</intersection>
<intersection>1363 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>454,1363,455,1363</points>
<connection>
<GID>1253</GID>
<name>IN_0</name></connection>
<intersection>454 4</intersection></hsegment></shape></wire>
<wire>
<ID>1864</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,1361,455,1361</points>
<connection>
<GID>1254</GID>
<name>IN_0</name></connection>
<intersection>454.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>454.5,1360,454.5,1361</points>
<intersection>1360 4</intersection>
<intersection>1361 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>449,1360,454.5,1360</points>
<connection>
<GID>1244</GID>
<name>OUT_1</name></connection>
<intersection>454.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>1865</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>449,1359,455,1359</points>
<connection>
<GID>1244</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1255</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1866</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>562.5,1382.5,562.5,1390.5</points>
<connection>
<GID>1256</GID>
<name>IN_0</name></connection>
<intersection>1390.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>562.5,1390.5,566.5,1390.5</points>
<connection>
<GID>1104</GID>
<name>IN_7</name></connection>
<intersection>562.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1867</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563,1380.5,563,1389.5</points>
<intersection>1380.5 2</intersection>
<intersection>1389.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>563,1389.5,566.5,1389.5</points>
<connection>
<GID>1104</GID>
<name>IN_6</name></connection>
<intersection>563 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>562.5,1380.5,563,1380.5</points>
<connection>
<GID>1257</GID>
<name>IN_0</name></connection>
<intersection>563 0</intersection></hsegment></shape></wire>
<wire>
<ID>1868</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>566,1368.5,566,1383.5</points>
<intersection>1368.5 1</intersection>
<intersection>1383.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1368.5,566,1368.5</points>
<connection>
<GID>1264</GID>
<name>IN_0</name></connection>
<intersection>566 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>566,1383.5,566.5,1383.5</points>
<connection>
<GID>1104</GID>
<name>IN_0</name></connection>
<intersection>566 0</intersection></hsegment></shape></wire>
<wire>
<ID>1869</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565.5,1370.5,565.5,1384.5</points>
<intersection>1370.5 1</intersection>
<intersection>1384.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1370.5,565.5,1370.5</points>
<connection>
<GID>1263</GID>
<name>IN_0</name></connection>
<intersection>565.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>565.5,1384.5,566.5,1384.5</points>
<connection>
<GID>1104</GID>
<name>IN_1</name></connection>
<intersection>565.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1870</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565,1372.5,565,1385.5</points>
<intersection>1372.5 1</intersection>
<intersection>1385.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1372.5,565,1372.5</points>
<connection>
<GID>1262</GID>
<name>IN_0</name></connection>
<intersection>565 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>565,1385.5,566.5,1385.5</points>
<connection>
<GID>1104</GID>
<name>IN_2</name></connection>
<intersection>565 0</intersection></hsegment></shape></wire>
<wire>
<ID>1871</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,1374.5,564.5,1386.5</points>
<intersection>1374.5 1</intersection>
<intersection>1386.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1374.5,564.5,1374.5</points>
<connection>
<GID>1260</GID>
<name>IN_0</name></connection>
<intersection>564.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>564.5,1386.5,566.5,1386.5</points>
<connection>
<GID>1104</GID>
<name>IN_3</name></connection>
<intersection>564.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1872</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564,1376.5,564,1387.5</points>
<intersection>1376.5 1</intersection>
<intersection>1387.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1376.5,564,1376.5</points>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection>
<intersection>564 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>564,1387.5,566.5,1387.5</points>
<connection>
<GID>1104</GID>
<name>IN_4</name></connection>
<intersection>564 0</intersection></hsegment></shape></wire>
<wire>
<ID>1873</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563.5,1378.5,563.5,1388.5</points>
<intersection>1378.5 1</intersection>
<intersection>1388.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>562.5,1378.5,563.5,1378.5</points>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection>
<intersection>563.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>563.5,1388.5,566.5,1388.5</points>
<connection>
<GID>1104</GID>
<name>IN_5</name></connection>
<intersection>563.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1874</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,1392.5,569.5,1395.5</points>
<connection>
<GID>1266</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1104</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>1875</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540,1327,540,1339</points>
<intersection>1327 1</intersection>
<intersection>1339 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1327,540,1327</points>
<connection>
<GID>1420</GID>
<name>OUT_4</name></connection>
<intersection>540 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540,1339,589.5,1339</points>
<connection>
<GID>1439</GID>
<name>IN_4</name></connection>
<intersection>540 0</intersection></hsegment></shape></wire>
<wire>
<ID>1876</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697.5,1378,697.5,1378</points>
<connection>
<GID>1268</GID>
<name>carry_out</name></connection>
<connection>
<GID>1269</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>1877</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1374.5,640.5,1374.5</points>
<connection>
<GID>1270</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1878</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>693.5,1372,694.5,1372</points>
<connection>
<GID>1269</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>1272</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1879</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>693.5,1373,693.5,1374</points>
<connection>
<GID>1273</GID>
<name>IN_0</name></connection>
<intersection>1373 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>693.5,1373,694.5,1373</points>
<connection>
<GID>1269</GID>
<name>IN_B_2</name></connection>
<intersection>693.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1880</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>693.5,1376,694,1376</points>
<connection>
<GID>1274</GID>
<name>IN_0</name></connection>
<intersection>694 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>694,1374,694,1376</points>
<intersection>1374 4</intersection>
<intersection>1376 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>694,1374,694.5,1374</points>
<connection>
<GID>1269</GID>
<name>IN_B_1</name></connection>
<intersection>694 3</intersection></hsegment></shape></wire>
<wire>
<ID>1881</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694.5,1375,694.5,1378</points>
<connection>
<GID>1269</GID>
<name>IN_B_0</name></connection>
<intersection>1378 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>693.5,1378,694.5,1378</points>
<connection>
<GID>1275</GID>
<name>IN_0</name></connection>
<intersection>694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1882</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>677.5,1371.5,677.5,1391</points>
<intersection>1371.5 2</intersection>
<intersection>1391 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>677.5,1391,694.5,1391</points>
<connection>
<GID>1268</GID>
<name>IN_B_0</name></connection>
<intersection>677.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638,1371.5,677.5,1371.5</points>
<connection>
<GID>1270</GID>
<name>OUT_0</name></connection>
<intersection>677.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1883</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>677,1372.5,677,1390</points>
<intersection>1372.5 2</intersection>
<intersection>1390 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>677,1390,694.5,1390</points>
<connection>
<GID>1268</GID>
<name>IN_B_1</name></connection>
<intersection>677 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638,1372.5,677,1372.5</points>
<connection>
<GID>1270</GID>
<name>OUT_1</name></connection>
<intersection>677 0</intersection></hsegment></shape></wire>
<wire>
<ID>1884</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>676.5,1373.5,676.5,1389</points>
<intersection>1373.5 2</intersection>
<intersection>1389 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>676.5,1389,694.5,1389</points>
<connection>
<GID>1268</GID>
<name>IN_B_2</name></connection>
<intersection>676.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>638,1373.5,676.5,1373.5</points>
<connection>
<GID>1270</GID>
<name>OUT_2</name></connection>
<intersection>676.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1885</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>693.5,1388,694.5,1388</points>
<connection>
<GID>1268</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>1276</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1886</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>693.5,1386,694.5,1386</points>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection>
<intersection>694.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>694.5,1384,694.5,1386</points>
<connection>
<GID>1268</GID>
<name>IN_0</name></connection>
<intersection>1386 7</intersection></vsegment></shape></wire>
<wire>
<ID>1887</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694,1383,694,1384</points>
<intersection>1383 5</intersection>
<intersection>1384 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>693.5,1384,694,1384</points>
<connection>
<GID>1283</GID>
<name>IN_0</name></connection>
<intersection>694 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>694,1383,694.5,1383</points>
<connection>
<GID>1268</GID>
<name>IN_1</name></connection>
<intersection>694 0</intersection></hsegment></shape></wire>
<wire>
<ID>1888</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>693.5,1382,694.5,1382</points>
<connection>
<GID>1268</GID>
<name>IN_2</name></connection>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1889</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694.5,1380,694.5,1381</points>
<connection>
<GID>1268</GID>
<name>IN_3</name></connection>
<intersection>1380 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>693.5,1380,694.5,1380</points>
<connection>
<GID>1282</GID>
<name>IN_0</name></connection>
<intersection>694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1890</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>693.5,1370,694.5,1370</points>
<connection>
<GID>1280</GID>
<name>IN_0</name></connection>
<intersection>694.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>694.5,1368,694.5,1370</points>
<connection>
<GID>1269</GID>
<name>IN_0</name></connection>
<intersection>1370 1</intersection></vsegment></shape></wire>
<wire>
<ID>1891</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694,1367,694,1368</points>
<intersection>1367 2</intersection>
<intersection>1368 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>693.5,1368,694,1368</points>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection>
<intersection>694 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>694,1367,694.5,1367</points>
<connection>
<GID>1269</GID>
<name>IN_1</name></connection>
<intersection>694 0</intersection></hsegment></shape></wire>
<wire>
<ID>1892</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>693.5,1366,694.5,1366</points>
<connection>
<GID>1269</GID>
<name>IN_2</name></connection>
<connection>
<GID>1278</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1893</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694.5,1364,694.5,1365</points>
<connection>
<GID>1269</GID>
<name>IN_3</name></connection>
<intersection>1364 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>693.5,1364,694.5,1364</points>
<connection>
<GID>1277</GID>
<name>IN_0</name></connection>
<intersection>694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1894</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539.5,1328,539.5,1340</points>
<intersection>1328 1</intersection>
<intersection>1340 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1328,539.5,1328</points>
<connection>
<GID>1420</GID>
<name>OUT_5</name></connection>
<intersection>539.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539.5,1340,589.5,1340</points>
<connection>
<GID>1439</GID>
<name>IN_5</name></connection>
<intersection>539.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1895</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>447,1367.5,447,1368.5</points>
<connection>
<GID>1244</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1248</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1896</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>702.5,1387.5,702.5,1389</points>
<connection>
<GID>1268</GID>
<name>OUT_0</name></connection>
<intersection>1389 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>702.5,1389,703,1389</points>
<connection>
<GID>1306</GID>
<name>IN_0</name></connection>
<intersection>702.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1897</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>702.5,1387,703,1387</points>
<connection>
<GID>1307</GID>
<name>IN_0</name></connection>
<intersection>702.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>702.5,1386.5,702.5,1387</points>
<connection>
<GID>1268</GID>
<name>OUT_1</name></connection>
<intersection>1387 0</intersection></vsegment></shape></wire>
<wire>
<ID>1898</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>702.5,1385,702.5,1385.5</points>
<connection>
<GID>1268</GID>
<name>OUT_2</name></connection>
<intersection>1385 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>702.5,1385,703,1385</points>
<connection>
<GID>1308</GID>
<name>IN_0</name></connection>
<intersection>702.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1899</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>702.5,1383,702.5,1384.5</points>
<connection>
<GID>1268</GID>
<name>OUT_3</name></connection>
<intersection>1383 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>702.5,1383,703,1383</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<intersection>702.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1900</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>702.5,1371.5,702.5,1373</points>
<connection>
<GID>1269</GID>
<name>OUT_0</name></connection>
<intersection>1373 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>702.5,1373,703,1373</points>
<connection>
<GID>1310</GID>
<name>IN_0</name></connection>
<intersection>702.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1901</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>702.5,1370.5,702.5,1371</points>
<connection>
<GID>1269</GID>
<name>OUT_1</name></connection>
<intersection>1371 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>702.5,1371,703,1371</points>
<connection>
<GID>1311</GID>
<name>IN_0</name></connection>
<intersection>702.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1902</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>702.5,1369,703,1369</points>
<connection>
<GID>1312</GID>
<name>IN_0</name></connection>
<intersection>702.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>702.5,1369,702.5,1369.5</points>
<connection>
<GID>1269</GID>
<name>OUT_2</name></connection>
<intersection>1369 8</intersection></vsegment></shape></wire>
<wire>
<ID>1903</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>702.5,1367,702.5,1368.5</points>
<connection>
<GID>1269</GID>
<name>OUT_3</name></connection>
<intersection>1367 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>702.5,1367,703,1367</points>
<connection>
<GID>1313</GID>
<name>IN_0</name></connection>
<intersection>702.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1904</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,1381,426.5,1388</points>
<intersection>1381 4</intersection>
<intersection>1388 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>426.5,1381,428,1381</points>
<connection>
<GID>1302</GID>
<name>IN_7</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>423,1388,426.5,1388</points>
<connection>
<GID>1317</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1905</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423,1386,426,1386</points>
<connection>
<GID>1319</GID>
<name>IN_0</name></connection>
<intersection>426 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>426,1380,426,1386</points>
<intersection>1380 7</intersection>
<intersection>1386 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>426,1380,428,1380</points>
<connection>
<GID>1302</GID>
<name>IN_6</name></connection>
<intersection>426 4</intersection></hsegment></shape></wire>
<wire>
<ID>1906</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1379,425.5,1384</points>
<intersection>1379 4</intersection>
<intersection>1384 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,1384,425.5,1384</points>
<connection>
<GID>1320</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>425.5,1379,428,1379</points>
<connection>
<GID>1302</GID>
<name>IN_5</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1907</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423,1382,425,1382</points>
<connection>
<GID>1321</GID>
<name>IN_0</name></connection>
<intersection>425 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>425,1378,425,1382</points>
<intersection>1378 7</intersection>
<intersection>1382 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>425,1378,428,1378</points>
<connection>
<GID>1302</GID>
<name>IN_4</name></connection>
<intersection>425 4</intersection></hsegment></shape></wire>
<wire>
<ID>1908</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>423,1380,424.5,1380</points>
<connection>
<GID>1322</GID>
<name>IN_0</name></connection>
<intersection>424.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>424.5,1377,424.5,1380</points>
<intersection>1377 11</intersection>
<intersection>1380 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>424.5,1377,428,1377</points>
<connection>
<GID>1302</GID>
<name>IN_3</name></connection>
<intersection>424.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>1909</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>424,1376,424,1378</points>
<intersection>1376 7</intersection>
<intersection>1378 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>424,1376,428,1376</points>
<connection>
<GID>1302</GID>
<name>IN_2</name></connection>
<intersection>424 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>423,1378,424,1378</points>
<connection>
<GID>1323</GID>
<name>IN_0</name></connection>
<intersection>424 4</intersection></hsegment></shape></wire>
<wire>
<ID>1910</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,1375,423.5,1376</points>
<intersection>1375 4</intersection>
<intersection>1376 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,1376,423.5,1376</points>
<connection>
<GID>1324</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>423.5,1375,428,1375</points>
<connection>
<GID>1302</GID>
<name>IN_1</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1911</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423,1374,428,1374</points>
<connection>
<GID>1302</GID>
<name>IN_0</name></connection>
<connection>
<GID>1325</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1912</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,1329,539,1341</points>
<intersection>1329 1</intersection>
<intersection>1341 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1329,539,1329</points>
<connection>
<GID>1420</GID>
<name>OUT_6</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,1341,589.5,1341</points>
<connection>
<GID>1439</GID>
<name>IN_6</name></connection>
<intersection>539 0</intersection></hsegment></shape></wire>
<wire>
<ID>1913</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>667.5,1404,667.5,1404</points>
<connection>
<GID>1328</GID>
<name>carry_out</name></connection>
<connection>
<GID>1329</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>1914</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,1326,540.5,1338</points>
<intersection>1326 1</intersection>
<intersection>1338 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1326,540.5,1326</points>
<connection>
<GID>1420</GID>
<name>OUT_3</name></connection>
<intersection>540.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>540.5,1338,589.5,1338</points>
<connection>
<GID>1439</GID>
<name>IN_3</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532,1342,532,1347</points>
<intersection>1342 2</intersection>
<intersection>1347 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>532,1347,558,1347</points>
<connection>
<GID>1015</GID>
<name>IN_2</name></connection>
<intersection>532 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,1342,532,1342</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<intersection>532 0</intersection></hsegment></shape></wire>
<wire>
<ID>1915</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541.5,1324,541.5,1336</points>
<intersection>1324 1</intersection>
<intersection>1336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1324,541.5,1324</points>
<connection>
<GID>1420</GID>
<name>OUT_1</name></connection>
<intersection>541.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541.5,1336,589.5,1336</points>
<connection>
<GID>1439</GID>
<name>IN_1</name></connection>
<intersection>541.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1916</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541,1325,541,1337</points>
<intersection>1325 1</intersection>
<intersection>1337 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>511,1325,541,1325</points>
<connection>
<GID>1420</GID>
<name>OUT_2</name></connection>
<intersection>541 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>541,1337,589.5,1337</points>
<connection>
<GID>1439</GID>
<name>IN_2</name></connection>
<intersection>541 0</intersection></hsegment></shape></wire>
<wire>
<ID>1917</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>590.5,1343.5,591.5,1343.5</points>
<connection>
<GID>1439</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1440</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1918</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1412.5,664.5,1414</points>
<connection>
<GID>1328</GID>
<name>IN_B_3</name></connection>
<intersection>1412.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1412.5,664.5,1412.5</points>
<connection>
<GID>1334</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1919</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1410,664.5,1410.5</points>
<connection>
<GID>1328</GID>
<name>IN_0</name></connection>
<intersection>1410.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1410.5,664.5,1410.5</points>
<connection>
<GID>1342</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532.5,1340,532.5,1346</points>
<intersection>1340 2</intersection>
<intersection>1346 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>532.5,1346,558,1346</points>
<connection>
<GID>1015</GID>
<name>IN_1</name></connection>
<intersection>532.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,1340,532.5,1340</points>
<connection>
<GID>1006</GID>
<name>IN_0</name></connection>
<intersection>532.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1920</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1408.5,664.5,1409</points>
<connection>
<GID>1328</GID>
<name>IN_1</name></connection>
<intersection>1408.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>664,1408.5,664.5,1408.5</points>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1921</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664,1406.5,664,1408</points>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection>
<intersection>1408 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>664,1408,664.5,1408</points>
<connection>
<GID>1328</GID>
<name>IN_2</name></connection>
<intersection>664 0</intersection></hsegment></shape></wire>
<wire>
<ID>1922</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1404.5,664.5,1407</points>
<connection>
<GID>1328</GID>
<name>IN_3</name></connection>
<intersection>1404.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>664,1404.5,664.5,1404.5</points>
<connection>
<GID>1340</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1923</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1394,664.5,1394.5</points>
<connection>
<GID>1329</GID>
<name>IN_0</name></connection>
<intersection>1394.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1394.5,664.5,1394.5</points>
<connection>
<GID>1338</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1924</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1392.5,664.5,1393</points>
<connection>
<GID>1329</GID>
<name>IN_1</name></connection>
<intersection>1392.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>664,1392.5,664.5,1392.5</points>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1925</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664,1390.5,664,1392</points>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection>
<intersection>1392 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>664,1392,664.5,1392</points>
<connection>
<GID>1329</GID>
<name>IN_2</name></connection>
<intersection>664 0</intersection></hsegment></shape></wire>
<wire>
<ID>1926</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1388.5,664.5,1391</points>
<connection>
<GID>1329</GID>
<name>IN_3</name></connection>
<intersection>1388.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>664,1388.5,664.5,1388.5</points>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1927</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672.5,1413.5,672.5,1415</points>
<connection>
<GID>1328</GID>
<name>OUT_0</name></connection>
<intersection>1415 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>672.5,1415,673,1415</points>
<connection>
<GID>1343</GID>
<name>IN_0</name></connection>
<intersection>672.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1928</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>672.5,1413,673,1413</points>
<connection>
<GID>1344</GID>
<name>IN_0</name></connection>
<intersection>672.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>672.5,1412.5,672.5,1413</points>
<connection>
<GID>1328</GID>
<name>OUT_1</name></connection>
<intersection>1413 1</intersection></vsegment></shape></wire>
<wire>
<ID>1929</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>672.5,1411,673,1411</points>
<connection>
<GID>1345</GID>
<name>IN_0</name></connection>
<intersection>672.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>672.5,1411,672.5,1411.5</points>
<connection>
<GID>1328</GID>
<name>OUT_2</name></connection>
<intersection>1411 1</intersection></vsegment></shape></wire>
<wire>
<ID>1930</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672.5,1409,672.5,1410.5</points>
<connection>
<GID>1328</GID>
<name>OUT_3</name></connection>
<intersection>1409 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>672.5,1409,673,1409</points>
<connection>
<GID>1346</GID>
<name>IN_0</name></connection>
<intersection>672.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1931</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672.5,1397.5,672.5,1399</points>
<connection>
<GID>1329</GID>
<name>OUT_0</name></connection>
<intersection>1399 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>672.5,1399,673,1399</points>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection>
<intersection>672.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1932</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>672.5,1397,673,1397</points>
<connection>
<GID>1348</GID>
<name>IN_0</name></connection>
<intersection>672.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>672.5,1396.5,672.5,1397</points>
<connection>
<GID>1329</GID>
<name>OUT_1</name></connection>
<intersection>1397 6</intersection></vsegment></shape></wire>
<wire>
<ID>1933</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>672.5,1395,673,1395</points>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection>
<intersection>672.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>672.5,1395,672.5,1395.5</points>
<connection>
<GID>1329</GID>
<name>OUT_2</name></connection>
<intersection>1395 0</intersection></vsegment></shape></wire>
<wire>
<ID>1934</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>672.5,1393,672.5,1394.5</points>
<connection>
<GID>1329</GID>
<name>OUT_3</name></connection>
<intersection>1393 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>672.5,1393,673,1393</points>
<connection>
<GID>1350</GID>
<name>IN_0</name></connection>
<intersection>672.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1935</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1401,664.5,1402.5</points>
<connection>
<GID>1329</GID>
<name>IN_B_0</name></connection>
<intersection>1402.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1402.5,664.5,1402.5</points>
<connection>
<GID>1351</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1936</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1400,664.5,1400.5</points>
<connection>
<GID>1329</GID>
<name>IN_B_1</name></connection>
<intersection>1400.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1400.5,664.5,1400.5</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1937</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1398.5,664.5,1399</points>
<connection>
<GID>1329</GID>
<name>IN_B_2</name></connection>
<intersection>1398.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>664,1398.5,664.5,1398.5</points>
<connection>
<GID>1353</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1938</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1396.5,664.5,1398</points>
<connection>
<GID>1329</GID>
<name>IN_B_3</name></connection>
<intersection>1396.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>664,1396.5,664.5,1396.5</points>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1939</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1414.5,664.5,1415</points>
<connection>
<GID>1328</GID>
<name>IN_B_2</name></connection>
<intersection>1414.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>664,1414.5,664.5,1414.5</points>
<connection>
<GID>1355</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1940</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>638.5,1390.5,638.5,1390.5</points>
<connection>
<GID>1326</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1356</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1941</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>650.5,1388.5,650.5,1417</points>
<intersection>1388.5 1</intersection>
<intersection>1417 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638.5,1388.5,650.5,1388.5</points>
<connection>
<GID>1326</GID>
<name>OUT_0</name></connection>
<intersection>650.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>650.5,1417,664.5,1417</points>
<connection>
<GID>1328</GID>
<name>IN_B_0</name></connection>
<intersection>650.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1942</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>651,1389.5,651,1416</points>
<intersection>1389.5 1</intersection>
<intersection>1416 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>638.5,1389.5,651,1389.5</points>
<connection>
<GID>1326</GID>
<name>OUT_1</name></connection>
<intersection>651 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>651,1416,664.5,1416</points>
<connection>
<GID>1328</GID>
<name>IN_B_1</name></connection>
<intersection>651 0</intersection></hsegment></shape></wire>
<wire>
<ID>1173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1305.5,680.5,1309.5</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<intersection>1305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1305.5,692,1305.5</points>
<connection>
<GID>990</GID>
<name>IN_5</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1943</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>632.5,1380,632.5,1400.5</points>
<intersection>1380 2</intersection>
<intersection>1400.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,1400.5,632.5,1400.5</points>
<connection>
<GID>1358</GID>
<name>OUT_0</name></connection>
<intersection>632.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>632.5,1380,636,1380</points>
<connection>
<GID>1270</GID>
<name>ENABLE_0</name></connection>
<intersection>632.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1944</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>636.5,1397,636.5,1401.5</points>
<connection>
<GID>1326</GID>
<name>ENABLE_0</name></connection>
<intersection>1401.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>631,1401.5,636.5,1401.5</points>
<connection>
<GID>1358</GID>
<name>OUT_1</name></connection>
<intersection>636.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1947</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>659,1333,659,1333</points>
<connection>
<GID>1053</GID>
<name>OUT</name></connection>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1948</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>625,1400.5,625,1400.5</points>
<connection>
<GID>1358</GID>
<name>IN_0</name></connection>
<connection>
<GID>1366</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1949</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>625,1403.5,625,1403.5</points>
<connection>
<GID>1358</GID>
<name>ENABLE</name></connection>
<connection>
<GID>1368</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1950</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>619,1402.5,619,1402.5</points>
<connection>
<GID>1368</GID>
<name>IN_1</name></connection>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1951</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>649,1353,649,1360.5</points>
<intersection>1353 8</intersection>
<intersection>1360.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>649,1360.5,657.5,1360.5</points>
<connection>
<GID>1055</GID>
<name>ENABLE</name></connection>
<intersection>649 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>647.5,1353,653,1353</points>
<connection>
<GID>1371</GID>
<name>IN_0</name></connection>
<connection>
<GID>1054</GID>
<name>OUT</name></connection>
<intersection>649 0</intersection></hsegment></shape></wire>
<wire>
<ID>1952</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>619,1404.5,619,1404.5</points>
<connection>
<GID>1368</GID>
<name>IN_0</name></connection>
<connection>
<GID>1373</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1954</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,1369.5,489,1373.5</points>
<intersection>1369.5 2</intersection>
<intersection>1373.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1373.5,489,1373.5</points>
<connection>
<GID>1377</GID>
<name>IN_0</name></connection>
<intersection>489 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>489,1369.5,489.5,1369.5</points>
<connection>
<GID>1376</GID>
<name>IN_7</name></connection>
<intersection>489 0</intersection></hsegment></shape></wire>
<wire>
<ID>1955</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1371.5,488.5,1371.5</points>
<connection>
<GID>1378</GID>
<name>IN_0</name></connection>
<intersection>488.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>488.5,1368.5,488.5,1371.5</points>
<intersection>1368.5 5</intersection>
<intersection>1371.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>488.5,1368.5,489.5,1368.5</points>
<connection>
<GID>1376</GID>
<name>IN_6</name></connection>
<intersection>488.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1956</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488,1367.5,488,1369.5</points>
<intersection>1367.5 2</intersection>
<intersection>1369.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1369.5,488,1369.5</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<intersection>488 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488,1367.5,489.5,1367.5</points>
<connection>
<GID>1376</GID>
<name>IN_5</name></connection>
<intersection>488 0</intersection></hsegment></shape></wire>
<wire>
<ID>1957</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1367.5,487.5,1367.5</points>
<connection>
<GID>1380</GID>
<name>IN_0</name></connection>
<intersection>487.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>487.5,1366.5,487.5,1367.5</points>
<intersection>1366.5 5</intersection>
<intersection>1367.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>487.5,1366.5,489.5,1366.5</points>
<connection>
<GID>1376</GID>
<name>IN_4</name></connection>
<intersection>487.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1958</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>481.5,1365.5,489.5,1365.5</points>
<connection>
<GID>1376</GID>
<name>IN_3</name></connection>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1959</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1363.5,487.5,1363.5</points>
<connection>
<GID>1382</GID>
<name>IN_0</name></connection>
<intersection>487.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>487.5,1363.5,487.5,1364.5</points>
<intersection>1363.5 1</intersection>
<intersection>1364.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>487.5,1364.5,489.5,1364.5</points>
<connection>
<GID>1376</GID>
<name>IN_2</name></connection>
<intersection>487.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1960</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488,1361.5,488,1363.5</points>
<intersection>1361.5 1</intersection>
<intersection>1363.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1361.5,488,1361.5</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<intersection>488 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488,1363.5,489.5,1363.5</points>
<connection>
<GID>1376</GID>
<name>IN_1</name></connection>
<intersection>488 0</intersection></hsegment></shape></wire>
<wire>
<ID>1961</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488.5,1359.5,488.5,1362.5</points>
<intersection>1359.5 1</intersection>
<intersection>1362.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1359.5,488.5,1359.5</points>
<connection>
<GID>1384</GID>
<name>IN_0</name></connection>
<intersection>488.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488.5,1362.5,489.5,1362.5</points>
<connection>
<GID>1376</GID>
<name>IN_0</name></connection>
<intersection>488.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1962</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1371,491.5,1371</points>
<connection>
<GID>1376</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1385</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1963</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,1382.5,430,1382.5</points>
<connection>
<GID>1302</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1386</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1964</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>629.5,1350,686.5,1350</points>
<connection>
<GID>1108</GID>
<name>OUT_5</name></connection>
<intersection>649.5 6</intersection>
<intersection>686.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>686.5,1322.5,686.5,1350</points>
<intersection>1322.5 5</intersection>
<intersection>1350 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>686.5,1322.5,734,1322.5</points>
<connection>
<GID>1022</GID>
<name>IN_0</name></connection>
<intersection>686.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>649.5,1350,649.5,1358.5</points>
<intersection>1350 1</intersection>
<intersection>1358.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>649.5,1358.5,657.5,1358.5</points>
<connection>
<GID>1055</GID>
<name>IN_1</name></connection>
<intersection>649.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1968</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>556.5,1384.5,556.5,1393.5</points>
<intersection>1384.5 5</intersection>
<intersection>1393.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>556.5,1393.5,557,1393.5</points>
<connection>
<GID>1232</GID>
<name>IN_0</name></connection>
<intersection>556.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>553,1384.5,556.5,1384.5</points>
<connection>
<GID>1102</GID>
<name>OUT_1</name></connection>
<intersection>556.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1969</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>629.5,1349,686,1349</points>
<connection>
<GID>1108</GID>
<name>OUT_4</name></connection>
<intersection>650 6</intersection>
<intersection>686 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>686,1322,686,1349</points>
<intersection>1322 5</intersection>
<intersection>1349 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>686,1322,733.5,1322</points>
<intersection>686 4</intersection>
<intersection>733.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>650,1349,650,1357.5</points>
<intersection>1349 1</intersection>
<intersection>1357.5 9</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>733.5,1318.5,733.5,1322</points>
<intersection>1318.5 8</intersection>
<intersection>1322 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>733.5,1318.5,734,1318.5</points>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection>
<intersection>733.5 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>650,1357.5,657.5,1357.5</points>
<connection>
<GID>1055</GID>
<name>IN_0</name></connection>
<intersection>650 6</intersection></hsegment></shape></wire>
<wire>
<ID>1970</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1348,574.5,1348</points>
<connection>
<GID>1126</GID>
<name>IN_3</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1971</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1346,574.5,1346</points>
<connection>
<GID>1126</GID>
<name>IN_1</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1972</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1351,574.5,1351</points>
<connection>
<GID>1126</GID>
<name>IN_6</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1973</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1349,574.5,1349</points>
<connection>
<GID>1126</GID>
<name>IN_4</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1974</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1345,574.5,1345</points>
<connection>
<GID>1126</GID>
<name>IN_0</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1313.5,680.5,1317.5</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<intersection>1313.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1313.5,692,1313.5</points>
<connection>
<GID>990</GID>
<name>IN_13</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1976</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>626,1327,626,1334</points>
<intersection>1327 1</intersection>
<intersection>1334 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>626,1327,629.5,1327</points>
<connection>
<GID>1409</GID>
<name>IN_0</name></connection>
<intersection>626 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>620,1334,626,1334</points>
<connection>
<GID>1405</GID>
<name>OUT_0</name></connection>
<intersection>626 0</intersection></hsegment></shape></wire>
<wire>
<ID>1977</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>626.5,1329,626.5,1335</points>
<intersection>1329 1</intersection>
<intersection>1335 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>626.5,1329,629.5,1329</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<intersection>626.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>620,1335,626.5,1335</points>
<connection>
<GID>1405</GID>
<name>OUT_1</name></connection>
<intersection>626.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1978</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627,1331,627,1336</points>
<intersection>1331 7</intersection>
<intersection>1336 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>627,1331,629.5,1331</points>
<connection>
<GID>1413</GID>
<name>IN_0</name></connection>
<intersection>627 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>620,1336,627,1336</points>
<connection>
<GID>1405</GID>
<name>OUT_2</name></connection>
<intersection>627 0</intersection></hsegment></shape></wire>
<wire>
<ID>1979</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>627.5,1333,627.5,1337</points>
<intersection>1333 7</intersection>
<intersection>1337 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>620,1337,627.5,1337</points>
<connection>
<GID>1405</GID>
<name>OUT_3</name></connection>
<intersection>627.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>627.5,1333,629.5,1333</points>
<connection>
<GID>1414</GID>
<name>IN_0</name></connection>
<intersection>627.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1980</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>628,1335,629.5,1335</points>
<connection>
<GID>1415</GID>
<name>IN_0</name></connection>
<intersection>628 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>628,1335,628,1338</points>
<intersection>1335 2</intersection>
<intersection>1338 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>620,1338,628,1338</points>
<connection>
<GID>1405</GID>
<name>OUT_4</name></connection>
<intersection>628 6</intersection></hsegment></shape></wire>
<wire>
<ID>1981</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628.5,1337,628.5,1339</points>
<intersection>1337 1</intersection>
<intersection>1339 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>628.5,1337,629.5,1337</points>
<connection>
<GID>1416</GID>
<name>IN_0</name></connection>
<intersection>628.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>620,1339,628.5,1339</points>
<connection>
<GID>1405</GID>
<name>OUT_5</name></connection>
<intersection>628.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1982</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>620,1340,629,1340</points>
<connection>
<GID>1405</GID>
<name>OUT_6</name></connection>
<intersection>629 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>629,1339,629,1340</points>
<intersection>1339 12</intersection>
<intersection>1340 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>629,1339,629.5,1339</points>
<connection>
<GID>1417</GID>
<name>IN_0</name></connection>
<intersection>629 5</intersection></hsegment></shape></wire>
<wire>
<ID>1983</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>620,1341,629.5,1341</points>
<connection>
<GID>1405</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1418</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1984</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,1267,398,1274</points>
<intersection>1267 1</intersection>
<intersection>1274 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>394.5,1267,398,1267</points>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection>
<intersection>398 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>398,1274,409,1274</points>
<connection>
<GID>1109</GID>
<name>IN_0</name></connection>
<intersection>398 0</intersection></hsegment></shape></wire>
<wire>
<ID>1985</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394.5,1281,409,1281</points>
<connection>
<GID>1109</GID>
<name>IN_7</name></connection>
<connection>
<GID>1430</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1986</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>394.5,1279,395,1279</points>
<connection>
<GID>1429</GID>
<name>IN_0</name></connection>
<intersection>395 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>395,1279,395,1280</points>
<intersection>1279 1</intersection>
<intersection>1280 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>395,1280,409,1280</points>
<connection>
<GID>1109</GID>
<name>IN_6</name></connection>
<intersection>395 3</intersection></hsegment></shape></wire>
<wire>
<ID>1987</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395.5,1277,395.5,1279</points>
<intersection>1277 2</intersection>
<intersection>1279 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>395.5,1279,409,1279</points>
<connection>
<GID>1109</GID>
<name>IN_5</name></connection>
<intersection>395.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394.5,1277,395.5,1277</points>
<connection>
<GID>1428</GID>
<name>IN_0</name></connection>
<intersection>395.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1988</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396,1275,396,1278</points>
<intersection>1275 4</intersection>
<intersection>1278 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>396,1278,409,1278</points>
<connection>
<GID>1109</GID>
<name>IN_4</name></connection>
<intersection>396 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>394.5,1275,396,1275</points>
<connection>
<GID>1427</GID>
<name>IN_0</name></connection>
<intersection>396 0</intersection></hsegment></shape></wire>
<wire>
<ID>1989</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>396.5,1273,396.5,1277</points>
<intersection>1273 3</intersection>
<intersection>1277 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>396.5,1277,409,1277</points>
<connection>
<GID>1109</GID>
<name>IN_3</name></connection>
<intersection>396.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>394.5,1273,396.5,1273</points>
<connection>
<GID>1426</GID>
<name>IN_0</name></connection>
<intersection>396.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1990</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397,1271,397,1276</points>
<intersection>1271 2</intersection>
<intersection>1276 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>397,1276,409,1276</points>
<connection>
<GID>1109</GID>
<name>IN_2</name></connection>
<intersection>397 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394.5,1271,397,1271</points>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection>
<intersection>397 0</intersection></hsegment></shape></wire>
<wire>
<ID>1991</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>397.5,1269,397.5,1275</points>
<intersection>1269 2</intersection>
<intersection>1275 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>397.5,1275,409,1275</points>
<connection>
<GID>1109</GID>
<name>IN_1</name></connection>
<intersection>397.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>394.5,1269,397.5,1269</points>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection>
<intersection>397.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1992</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1347,574.5,1347</points>
<connection>
<GID>1126</GID>
<name>IN_2</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1993</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1350,574.5,1350</points>
<connection>
<GID>1126</GID>
<name>IN_5</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1994</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>562,1352,574.5,1352</points>
<connection>
<GID>1126</GID>
<name>IN_7</name></connection>
<connection>
<GID>1015</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1995</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>560,1353.5,560,1354</points>
<connection>
<GID>1015</GID>
<name>ENABLE_0</name></connection>
<intersection>1354 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>555,1354,560,1354</points>
<connection>
<GID>1454</GID>
<name>IN_0</name></connection>
<intersection>560 0</intersection></hsegment></shape></wire>
<wire>
<ID>1996</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>424.5,1312.5,427,1312.5</points>
<connection>
<GID>1298</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1997</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>706.5,1331,707,1331</points>
<connection>
<GID>1359</GID>
<name>IN_0</name></connection>
<intersection>706.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>706.5,1331,706.5,1332.5</points>
<connection>
<GID>1179</GID>
<name>OUT_3</name></connection>
<intersection>1331 1</intersection></vsegment></shape></wire>
<wire>
<ID>1998</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>697,1355,698.5,1355</points>
<connection>
<GID>1177</GID>
<name>IN_B_0</name></connection>
<intersection>697 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>697,1355,697,1355.5</points>
<connection>
<GID>1361</GID>
<name>OUT_0</name></connection>
<intersection>1355 4</intersection></vsegment></shape></wire>
<wire>
<ID>1999</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488.5,1386.5,488.5,1389.5</points>
<intersection>1386.5 2</intersection>
<intersection>1389.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1389.5,488.5,1389.5</points>
<connection>
<GID>1363</GID>
<name>IN_0</name></connection>
<intersection>488.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488.5,1386.5,489.5,1386.5</points>
<connection>
<GID>1362</GID>
<name>IN_7</name></connection>
<intersection>488.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2000</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1387.5,488,1387.5</points>
<connection>
<GID>1365</GID>
<name>IN_0</name></connection>
<intersection>488 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>488,1385.5,488,1387.5</points>
<intersection>1385.5 5</intersection>
<intersection>1387.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>488,1385.5,489.5,1385.5</points>
<connection>
<GID>1362</GID>
<name>IN_6</name></connection>
<intersection>488 4</intersection></hsegment></shape></wire>
<wire>
<ID>2001</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>401.5,1332,404,1332</points>
<connection>
<GID>1295</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2002</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411,1282.5,411,1285</points>
<connection>
<GID>1109</GID>
<name>ENABLE_0</name></connection>
<intersection>1285 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>409.5,1285,411,1285</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<intersection>411 0</intersection></hsegment></shape></wire>
<wire>
<ID>2003</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,1270,413.5,1270.5</points>
<connection>
<GID>1469</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1471</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2007</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1385.5,487.5,1385.5</points>
<connection>
<GID>1367</GID>
<name>IN_0</name></connection>
<intersection>487.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>487.5,1384.5,487.5,1385.5</points>
<intersection>1384.5 3</intersection>
<intersection>1385.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>487.5,1384.5,489.5,1384.5</points>
<connection>
<GID>1362</GID>
<name>IN_5</name></connection>
<intersection>487.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>2008</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1383.5,489.5,1383.5</points>
<connection>
<GID>1362</GID>
<name>IN_4</name></connection>
<connection>
<GID>1370</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2014</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>481.5,1381.5,487.5,1381.5</points>
<connection>
<GID>1372</GID>
<name>IN_0</name></connection>
<intersection>487.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>487.5,1381.5,487.5,1382.5</points>
<intersection>1381.5 7</intersection>
<intersection>1382.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>487.5,1382.5,489.5,1382.5</points>
<connection>
<GID>1362</GID>
<name>IN_3</name></connection>
<intersection>487.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>2015</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>406,1268.5,411.5,1268.5</points>
<connection>
<GID>1469</GID>
<name>IN_7</name></connection>
<connection>
<GID>1492</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2016</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>406.5,1266.5,406.5,1267.5</points>
<intersection>1266.5 1</intersection>
<intersection>1267.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1266.5,406.5,1266.5</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>406.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>406.5,1267.5,411.5,1267.5</points>
<connection>
<GID>1469</GID>
<name>IN_6</name></connection>
<intersection>406.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2017</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,1264.5,407,1266.5</points>
<intersection>1264.5 3</intersection>
<intersection>1266.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>407,1266.5,411.5,1266.5</points>
<connection>
<GID>1469</GID>
<name>IN_5</name></connection>
<intersection>407 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>406,1264.5,407,1264.5</points>
<connection>
<GID>1490</GID>
<name>IN_0</name></connection>
<intersection>407 0</intersection></hsegment></shape></wire>
<wire>
<ID>2018</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407.5,1262.5,407.5,1265.5</points>
<intersection>1262.5 1</intersection>
<intersection>1265.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1262.5,407.5,1262.5</points>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection>
<intersection>407.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>407.5,1265.5,411.5,1265.5</points>
<connection>
<GID>1469</GID>
<name>IN_4</name></connection>
<intersection>407.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2019</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408,1260.5,408,1264.5</points>
<intersection>1260.5 1</intersection>
<intersection>1264.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1260.5,408,1260.5</points>
<connection>
<GID>1488</GID>
<name>IN_0</name></connection>
<intersection>408 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>408,1264.5,411.5,1264.5</points>
<connection>
<GID>1469</GID>
<name>IN_3</name></connection>
<intersection>408 0</intersection></hsegment></shape></wire>
<wire>
<ID>2020</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,1258.5,408.5,1263.5</points>
<intersection>1258.5 1</intersection>
<intersection>1263.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1258.5,408.5,1258.5</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>408.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>408.5,1263.5,411.5,1263.5</points>
<connection>
<GID>1469</GID>
<name>IN_2</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>409,1256.5,409,1262.5</points>
<intersection>1256.5 1</intersection>
<intersection>1262.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1256.5,409,1256.5</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>409 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>409,1262.5,411.5,1262.5</points>
<connection>
<GID>1469</GID>
<name>IN_1</name></connection>
<intersection>409 0</intersection></hsegment></shape></wire>
<wire>
<ID>2022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>409.5,1254.5,409.5,1261.5</points>
<intersection>1254.5 1</intersection>
<intersection>1261.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>406,1254.5,409.5,1254.5</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<intersection>409.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>409.5,1261.5,411.5,1261.5</points>
<connection>
<GID>1469</GID>
<name>IN_0</name></connection>
<intersection>409.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2023</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>573.5,1331.5,576,1331.5</points>
<connection>
<GID>1496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1207</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>2024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411,1301,411,1320</points>
<intersection>1301 3</intersection>
<intersection>1320 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>411,1301,427.5,1301</points>
<connection>
<GID>1506</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1500</GID>
<name>OUT</name></connection>
<intersection>411 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>404,1320,411,1320</points>
<connection>
<GID>1498</GID>
<name>ENABLE_0</name></connection>
<intersection>411 0</intersection></hsegment></shape></wire>
<wire>
<ID>2025</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>405,1302,405,1302</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2026</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>405,1300,405,1300</points>
<connection>
<GID>1500</GID>
<name>IN_1</name></connection>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1297.5,425.5,1298</points>
<connection>
<GID>1506</GID>
<name>IN_1</name></connection>
<intersection>1298 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424,1298,425.5,1298</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,1296,425.5,1296.5</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>1296 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424,1296,425.5,1296</points>
<connection>
<GID>1508</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2029</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>399.5,1318.5,402,1318.5</points>
<connection>
<GID>1498</GID>
<name>IN_3</name></connection>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400,1316.5,400,1317.5</points>
<intersection>1316.5 2</intersection>
<intersection>1317.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>400,1317.5,402,1317.5</points>
<connection>
<GID>1498</GID>
<name>IN_2</name></connection>
<intersection>400 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399.5,1316.5,400,1316.5</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>400 0</intersection></hsegment></shape></wire>
<wire>
<ID>2031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,1314.5,400.5,1316.5</points>
<intersection>1314.5 4</intersection>
<intersection>1316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>400.5,1316.5,402,1316.5</points>
<connection>
<GID>1498</GID>
<name>IN_1</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>399.5,1314.5,400.5,1314.5</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>400.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>401,1312.5,401,1315.5</points>
<intersection>1312.5 4</intersection>
<intersection>1315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>401,1315.5,402,1315.5</points>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection>
<intersection>401 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>399.5,1312.5,401,1312.5</points>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection>
<intersection>401 0</intersection></hsegment></shape></wire>
<wire>
<ID>2033</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1283,693,1283</points>
<connection>
<GID>1513</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>688 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>688,1283,688,1294</points>
<intersection>1283 1</intersection>
<intersection>1294 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>688,1294,711.5,1294</points>
<connection>
<GID>1075</GID>
<name>IN_1</name></connection>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection>
<intersection>688 7</intersection>
<intersection>699.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>699.5,1294,699.5,1315.5</points>
<intersection>1294 8</intersection>
<intersection>1315.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>696,1315.5,699.5,1315.5</points>
<connection>
<GID>990</GID>
<name>OUT_15</name></connection>
<intersection>699.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>2034</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1281,693,1281</points>
<connection>
<GID>1513</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>689 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>689,1281,689,1292</points>
<intersection>1281 1</intersection>
<intersection>1292 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>689,1292,704,1292</points>
<connection>
<GID>1060</GID>
<name>IN_2</name></connection>
<intersection>689 10</intersection>
<intersection>698.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>698.5,1292,698.5,1311.5</points>
<intersection>1292 11</intersection>
<intersection>1311.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>696,1311.5,698.5,1311.5</points>
<connection>
<GID>990</GID>
<name>OUT_11</name></connection>
<intersection>698.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>2035</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1279,693,1279</points>
<connection>
<GID>1513</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>690 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>690,1279,690,1290</points>
<intersection>1279 1</intersection>
<intersection>1290 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>690,1290,704,1290</points>
<connection>
<GID>1060</GID>
<name>IN_7</name></connection>
<intersection>690 7</intersection>
<intersection>697.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>697.5,1290,697.5,1307.5</points>
<intersection>1290 8</intersection>
<intersection>1307.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>696,1307.5,697.5,1307.5</points>
<connection>
<GID>990</GID>
<name>OUT_7</name></connection>
<intersection>697.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>2036</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1282,701,1282</points>
<connection>
<GID>1513</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>688.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>688.5,1282,688.5,1293</points>
<intersection>1282 1</intersection>
<intersection>1293 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>688.5,1293,704,1293</points>
<connection>
<GID>1060</GID>
<name>IN_1</name></connection>
<intersection>688.5 7</intersection>
<intersection>699 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>699,1293,699,1313.5</points>
<intersection>1293 8</intersection>
<intersection>1313.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>696,1313.5,699,1313.5</points>
<connection>
<GID>990</GID>
<name>OUT_13</name></connection>
<intersection>699 12</intersection></hsegment></shape></wire>
<wire>
<ID>2037</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1280,701,1280</points>
<connection>
<GID>1513</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection>
<intersection>689.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>689.5,1280,689.5,1291</points>
<intersection>1280 1</intersection>
<intersection>1291 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>689.5,1291,704,1291</points>
<connection>
<GID>1060</GID>
<name>IN_3</name></connection>
<intersection>689.5 7</intersection>
<intersection>698 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>698,1291,698,1309.5</points>
<intersection>1291 8</intersection>
<intersection>1309.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>696,1309.5,698,1309.5</points>
<connection>
<GID>990</GID>
<name>OUT_9</name></connection>
<intersection>698 12</intersection></hsegment></shape></wire>
<wire>
<ID>2038</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1278,701,1278</points>
<connection>
<GID>1513</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>690.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>690.5,1278,690.5,1289</points>
<intersection>1278 1</intersection>
<intersection>1289 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>690.5,1289,704,1289</points>
<connection>
<GID>1060</GID>
<name>IN_6</name></connection>
<intersection>690.5 7</intersection>
<intersection>697 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>697,1289,697,1305.5</points>
<intersection>1289 8</intersection>
<intersection>1305.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>696,1305.5,697,1305.5</points>
<connection>
<GID>990</GID>
<name>OUT_5</name></connection>
<intersection>697 12</intersection></hsegment></shape></wire>
<wire>
<ID>2039</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1277,693,1277</points>
<connection>
<GID>1513</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>691 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>691,1277,691,1288</points>
<intersection>1277 1</intersection>
<intersection>1288 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>691,1288,704,1288</points>
<connection>
<GID>1060</GID>
<name>IN_5</name></connection>
<intersection>691 10</intersection>
<intersection>696.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>696.5,1288,696.5,1303.5</points>
<intersection>1288 11</intersection>
<intersection>1303.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>696,1303.5,696.5,1303.5</points>
<connection>
<GID>990</GID>
<name>OUT_3</name></connection>
<intersection>696.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>2040</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673.5,1276,701,1276</points>
<connection>
<GID>1513</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>691.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>691.5,1276,691.5,1287</points>
<intersection>1276 1</intersection>
<intersection>1287 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>691.5,1287,704,1287</points>
<connection>
<GID>1060</GID>
<name>IN_4</name></connection>
<intersection>691.5 7</intersection>
<intersection>696 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>696,1287,696,1301.5</points>
<connection>
<GID>990</GID>
<name>OUT_1</name></connection>
<intersection>1287 12</intersection></vsegment></shape></wire>
<wire>
<ID>2041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>702,1284.5,702,1306.5</points>
<intersection>1284.5 3</intersection>
<intersection>1306.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>702,1306.5,726.5,1306.5</points>
<intersection>702 0</intersection>
<intersection>726.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>726.5,1305.5,726.5,1306.5</points>
<connection>
<GID>1549</GID>
<name>IN_0</name></connection>
<intersection>1306.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>671.5,1284.5,702,1284.5</points>
<connection>
<GID>1513</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1525</GID>
<name>OUT</name></connection>
<intersection>702 0</intersection></hsegment></shape></wire>
<wire>
<ID>2042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672.5,1290.5,672.5,1290.5</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>670.5,1290.5,670.5,1290.5</points>
<connection>
<GID>1525</GID>
<name>IN_1</name></connection>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2044</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>481.5,1379.5,488,1379.5</points>
<connection>
<GID>1374</GID>
<name>IN_0</name></connection>
<intersection>488 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>488,1379.5,488,1381.5</points>
<intersection>1379.5 1</intersection>
<intersection>1381.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>488,1381.5,489.5,1381.5</points>
<connection>
<GID>1362</GID>
<name>IN_2</name></connection>
<intersection>488 4</intersection></hsegment></shape></wire>
<wire>
<ID>2045</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>488.5,1377.5,488.5,1380.5</points>
<intersection>1377.5 1</intersection>
<intersection>1380.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1377.5,488.5,1377.5</points>
<connection>
<GID>1375</GID>
<name>IN_0</name></connection>
<intersection>488.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>488.5,1380.5,489.5,1380.5</points>
<connection>
<GID>1362</GID>
<name>IN_1</name></connection>
<intersection>488.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,1375.5,489,1379.5</points>
<intersection>1375.5 1</intersection>
<intersection>1379.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,1375.5,489,1375.5</points>
<connection>
<GID>1387</GID>
<name>IN_0</name></connection>
<intersection>489 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>489,1379.5,489.5,1379.5</points>
<connection>
<GID>1362</GID>
<name>IN_0</name></connection>
<intersection>489 0</intersection></hsegment></shape></wire>
<wire>
<ID>2052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1392,491.5,1392</points>
<connection>
<GID>1406</GID>
<name>IN_0</name></connection>
<connection>
<GID>1411</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2053</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1381.5,519,1381.5</points>
<connection>
<GID>1063</GID>
<name>IN_2</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_2</name></connection>
<intersection>496.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>496.5,1364.5,496.5,1381.5</points>
<intersection>1364.5 5</intersection>
<intersection>1381.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1364.5,496.5,1364.5</points>
<connection>
<GID>1376</GID>
<name>OUT_2</name></connection>
<intersection>496.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2054</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1383.5,519,1383.5</points>
<connection>
<GID>1362</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1063</GID>
<name>IN_4</name></connection>
<intersection>495.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>495.5,1366.5,495.5,1383.5</points>
<intersection>1366.5 5</intersection>
<intersection>1383.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1366.5,495.5,1366.5</points>
<connection>
<GID>1376</GID>
<name>OUT_4</name></connection>
<intersection>495.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2055</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1379.5,519,1379.5</points>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_0</name></connection>
<intersection>497.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>497.5,1362.5,497.5,1379.5</points>
<intersection>1362.5 5</intersection>
<intersection>1379.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1362.5,497.5,1362.5</points>
<connection>
<GID>1376</GID>
<name>OUT_0</name></connection>
<intersection>497.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2056</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1384.5,519,1384.5</points>
<connection>
<GID>1063</GID>
<name>IN_5</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_5</name></connection>
<intersection>495 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>495,1367.5,495,1384.5</points>
<intersection>1367.5 5</intersection>
<intersection>1384.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1367.5,495,1367.5</points>
<connection>
<GID>1376</GID>
<name>OUT_5</name></connection>
<intersection>495 4</intersection></hsegment></shape></wire>
<wire>
<ID>2057</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1380.5,519,1380.5</points>
<connection>
<GID>1063</GID>
<name>IN_1</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_1</name></connection>
<intersection>497 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>497,1363.5,497,1380.5</points>
<intersection>1363.5 5</intersection>
<intersection>1380.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1363.5,497,1363.5</points>
<connection>
<GID>1376</GID>
<name>OUT_1</name></connection>
<intersection>497 4</intersection></hsegment></shape></wire>
<wire>
<ID>2058</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1382.5,519,1382.5</points>
<connection>
<GID>1063</GID>
<name>IN_3</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_3</name></connection>
<intersection>496 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>496,1365.5,496,1382.5</points>
<intersection>1365.5 5</intersection>
<intersection>1382.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1365.5,496,1365.5</points>
<connection>
<GID>1376</GID>
<name>OUT_3</name></connection>
<intersection>496 4</intersection></hsegment></shape></wire>
<wire>
<ID>2059</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1385.5,519,1385.5</points>
<connection>
<GID>1063</GID>
<name>IN_6</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_6</name></connection>
<intersection>494.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>494.5,1368.5,494.5,1385.5</points>
<intersection>1368.5 5</intersection>
<intersection>1385.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1368.5,494.5,1368.5</points>
<connection>
<GID>1376</GID>
<name>OUT_6</name></connection>
<intersection>494.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>2060</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493.5,1386.5,519,1386.5</points>
<connection>
<GID>1063</GID>
<name>IN_7</name></connection>
<connection>
<GID>1362</GID>
<name>OUT_7</name></connection>
<intersection>494 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>494,1369.5,494,1386.5</points>
<intersection>1369.5 5</intersection>
<intersection>1386.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>493.5,1369.5,494,1369.5</points>
<connection>
<GID>1376</GID>
<name>OUT_7</name></connection>
<intersection>494 4</intersection></hsegment></shape></wire>
<wire>
<ID>2062</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1352,621.5,1352</points>
<connection>
<GID>1108</GID>
<name>IN_7</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>2063</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1349,621.5,1349</points>
<connection>
<GID>1108</GID>
<name>IN_4</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>2064</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1345,621.5,1345</points>
<connection>
<GID>1108</GID>
<name>IN_0</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2065</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1348,621.5,1348</points>
<connection>
<GID>1108</GID>
<name>IN_3</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>2066</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1350,621.5,1350</points>
<connection>
<GID>1108</GID>
<name>IN_5</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>2067</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1347,621.5,1347</points>
<connection>
<GID>1108</GID>
<name>IN_2</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>2068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1346,621.5,1346</points>
<connection>
<GID>1108</GID>
<name>IN_1</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>2069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619.5,1351,621.5,1351</points>
<connection>
<GID>1108</GID>
<name>IN_6</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>2070</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,1342.5,407,1342.5</points>
<connection>
<GID>1532</GID>
<name>IN_0</name></connection>
<intersection>1342.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407,1342.5,407,1342.5</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>407 0</intersection></hsegment></shape></wire>
<wire>
<ID>2071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,1340.5,407,1340.5</points>
<connection>
<GID>1532</GID>
<name>IN_1</name></connection>
<intersection>1340.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407,1340.5,407,1340.5</points>
<connection>
<GID>1536</GID>
<name>IN_0</name></connection>
<intersection>407 0</intersection></hsegment></shape></wire>
<wire>
<ID>2072</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607,1354,607,1354</points>
<connection>
<GID>1106</GID>
<name>load</name></connection>
<connection>
<GID>1438</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407,1338.5,407,1338.5</points>
<connection>
<GID>1532</GID>
<name>IN_2</name></connection>
<intersection>1338.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407,1338.5,407,1338.5</points>
<connection>
<GID>1538</GID>
<name>IN_0</name></connection>
<intersection>407 0</intersection></hsegment></shape></wire>
<wire>
<ID>2074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413,1340.5,413,1340.5</points>
<connection>
<GID>1532</GID>
<name>OUT</name></connection>
<intersection>1340.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413,1340.5,413,1340.5</points>
<connection>
<GID>1540</GID>
<name>IN_0</name></connection>
<intersection>413 0</intersection></hsegment></shape></wire>
<wire>
<ID>2075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548,1374,548,1381.5</points>
<connection>
<GID>1102</GID>
<name>clock</name></connection>
<intersection>1374 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>546.5,1374,548,1374</points>
<connection>
<GID>1129</GID>
<name>OUT</name></connection>
<intersection>548 0</intersection></hsegment></shape></wire>
<wire>
<ID>2076</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>428.5,1371.5,430,1371.5</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<connection>
<GID>1541</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2077</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,1388,491.5,1388</points>
<connection>
<GID>1362</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1406</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2078</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,1355.5,423.5,1360.5</points>
<intersection>1355.5 2</intersection>
<intersection>1360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423.5,1360.5,428,1360.5</points>
<connection>
<GID>1235</GID>
<name>IN_2</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421,1355.5,423.5,1355.5</points>
<connection>
<GID>1240</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423,1357.5,423,1361.5</points>
<intersection>1357.5 2</intersection>
<intersection>1361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423,1361.5,428,1361.5</points>
<connection>
<GID>1235</GID>
<name>IN_3</name></connection>
<intersection>423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421,1357.5,423,1357.5</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<intersection>423 0</intersection></hsegment></shape></wire>
<wire>
<ID>2080</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>548,1392.5,548,1392.5</points>
<connection>
<GID>1102</GID>
<name>load</name></connection>
<connection>
<GID>1547</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2082</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>534,1313,570.5,1313</points>
<connection>
<GID>1289</GID>
<name>IN_7</name></connection>
<connection>
<GID>1192</GID>
<name>OUT_3</name></connection>
<intersection>565 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>565,1290,565,1313</points>
<intersection>1290 4</intersection>
<intersection>1313 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>565,1290,570.5,1290</points>
<connection>
<GID>1290</GID>
<name>IN_7</name></connection>
<intersection>565 3</intersection></hsegment></shape></wire>
<wire>
<ID>2083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>536,1314,536,1315</points>
<intersection>1314 2</intersection>
<intersection>1315 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>536,1315,570.5,1315</points>
<connection>
<GID>1289</GID>
<name>IN_9</name></connection>
<intersection>536 0</intersection>
<intersection>564 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,1314,536,1314</points>
<connection>
<GID>1192</GID>
<name>OUT_4</name></connection>
<intersection>536 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>564,1292,564,1315</points>
<intersection>1292 4</intersection>
<intersection>1315 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>564,1292,570.5,1292</points>
<connection>
<GID>1290</GID>
<name>IN_9</name></connection>
<intersection>564 3</intersection></hsegment></shape></wire>
<wire>
<ID>2084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535.5,1315,535.5,1317</points>
<intersection>1315 2</intersection>
<intersection>1317 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535.5,1317,570.5,1317</points>
<connection>
<GID>1289</GID>
<name>IN_11</name></connection>
<intersection>535.5 0</intersection>
<intersection>563 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,1315,535.5,1315</points>
<connection>
<GID>1192</GID>
<name>OUT_5</name></connection>
<intersection>535.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>563,1294,563,1317</points>
<intersection>1294 4</intersection>
<intersection>1317 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>563,1294,570.5,1294</points>
<connection>
<GID>1290</GID>
<name>IN_11</name></connection>
<intersection>563 3</intersection></hsegment></shape></wire>
<wire>
<ID>2085</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535,1316,535,1319</points>
<intersection>1316 2</intersection>
<intersection>1319 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535,1319,570.5,1319</points>
<connection>
<GID>1289</GID>
<name>IN_13</name></connection>
<intersection>535 0</intersection>
<intersection>562 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,1316,535,1316</points>
<connection>
<GID>1192</GID>
<name>OUT_6</name></connection>
<intersection>535 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>562,1296,562,1319</points>
<intersection>1296 4</intersection>
<intersection>1319 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>562,1296,570.5,1296</points>
<connection>
<GID>1290</GID>
<name>IN_13</name></connection>
<intersection>562 3</intersection></hsegment></shape></wire>
<wire>
<ID>2086</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,1342.5,618,1342.5</points>
<connection>
<GID>1405</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1479</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2087</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617.5,1353.5,617.5,1353.5</points>
<connection>
<GID>1422</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1481</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2088</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>624.5,1354,624.5,1355.5</points>
<connection>
<GID>1108</GID>
<name>load</name></connection>
<intersection>1355.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>624,1355.5,624.5,1355.5</points>
<connection>
<GID>1483</GID>
<name>OUT_0</name></connection>
<intersection>624.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2089</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534.5,1317,534.5,1321</points>
<intersection>1317 2</intersection>
<intersection>1321 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534.5,1321,570.5,1321</points>
<connection>
<GID>1289</GID>
<name>IN_15</name></connection>
<intersection>534.5 0</intersection>
<intersection>561 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,1317,534.5,1317</points>
<connection>
<GID>1192</GID>
<name>OUT_7</name></connection>
<intersection>534.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>561,1298,561,1321</points>
<intersection>1298 4</intersection>
<intersection>1321 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>561,1298,570.5,1298</points>
<connection>
<GID>1290</GID>
<name>IN_15</name></connection>
<intersection>561 3</intersection></hsegment></shape></wire>
<wire>
<ID>2090</ID>
<shape>
<vsegment>
<ID>15</ID>
<points>430,1367,430,1367.5</points>
<connection>
<GID>1235</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1493</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2091</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>725.5,1299,725.5,1299.5</points>
<connection>
<GID>1084</GID>
<name>load</name></connection>
<connection>
<GID>1549</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>2092</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>663.5,1358,665,1358</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<intersection>663.5 3</intersection>
<intersection>664 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>663.5,1358,663.5,1358.5</points>
<connection>
<GID>1055</GID>
<name>OUT_1</name></connection>
<intersection>1358 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>664,1352.5,664,1358</points>
<intersection>1352.5 5</intersection>
<intersection>1358 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>664,1352.5,665.5,1352.5</points>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection>
<intersection>664 4</intersection></hsegment></shape></wire>
<wire>
<ID>2093</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>663.5,1360.5,663.5,1362</points>
<connection>
<GID>1055</GID>
<name>OUT_3</name></connection>
<intersection>1362 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>663.5,1362,665,1362</points>
<connection>
<GID>847</GID>
<name>IN_0</name></connection>
<intersection>663.5 0</intersection>
<intersection>664 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>664,1362,664,1365.5</points>
<intersection>1362 1</intersection>
<intersection>1365.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>664,1365.5,665.5,1365.5</points>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection>
<intersection>664 2</intersection></hsegment></shape></wire>
<wire>
<ID>2094</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402,1327.5,402,1327.5</points>
<connection>
<GID>1295</GID>
<name>IN_0</name></connection>
<intersection>1327.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402,1327.5,402,1327.5</points>
<connection>
<GID>1555</GID>
<name>IN_0</name></connection>
<intersection>402 0</intersection></hsegment></shape></wire>
<wire>
<ID>2095</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425,1308,425,1308</points>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection>
<intersection>1308 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425,1308,425,1308</points>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection>
<intersection>425 0</intersection></hsegment></shape></wire>
<wire>
<ID>2096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,1373,540.5,1373</points>
<connection>
<GID>1129</GID>
<name>IN_1</name></connection>
<intersection>1373 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540.5,1373,540.5,1373</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,1381.5,569.5,1381.5</points>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection>
<intersection>1381.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569.5,1381.5,569.5,1381.5</points>
<connection>
<GID>1104</GID>
<name>clock</name></connection>
<intersection>569.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2098</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>590,1388.5,590,1388.5</points>
<connection>
<GID>1107</GID>
<name>write_clock</name></connection>
<intersection>1388.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>590,1388.5,590,1388.5</points>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection>
<intersection>590 0</intersection></hsegment></shape></wire>
<wire>
<ID>2099</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>607,1343,624.5,1343</points>
<connection>
<GID>1108</GID>
<name>clock</name></connection>
<connection>
<GID>1106</GID>
<name>clock</name></connection>
<intersection>607 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>607,1342,607,1343</points>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection>
<intersection>1343 3</intersection></vsegment></shape></wire>
<wire>
<ID>2100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>725.5,1288.5,725.5,1290</points>
<connection>
<GID>1084</GID>
<name>clock</name></connection>
<intersection>1288.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>725,1288.5,725.5,1288.5</points>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection>
<intersection>725.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534,1392,534,1393</points>
<connection>
<GID>1065</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1573</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680.5,1301.5,680.5,1305.5</points>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>1301.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>680.5,1301.5,692,1301.5</points>
<connection>
<GID>990</GID>
<name>IN_1</name></connection>
<intersection>680.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694,1317,694,1317.5</points>
<connection>
<GID>990</GID>
<name>ENABLE_0</name></connection>
<intersection>1317.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>691.5,1317.5,724.5,1317.5</points>
<connection>
<GID>993</GID>
<name>IN_0</name></connection>
<intersection>694 0</intersection>
<intersection>724.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>724.5,1305.5,724.5,1317.5</points>
<connection>
<GID>1549</GID>
<name>IN_1</name></connection>
<intersection>1317.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>740,1313.5,740,1315.5</points>
<connection>
<GID>1028</GID>
<name>OUT</name></connection>
<intersection>1315.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>740,1315.5,740.5,1315.5</points>
<connection>
<GID>1033</GID>
<name>IN_2</name></connection>
<intersection>740 0</intersection></hsegment></shape></wire>
<wire>
<ID>1493</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>740,1317.5,740.5,1317.5</points>
<connection>
<GID>1026</GID>
<name>OUT</name></connection>
<connection>
<GID>1033</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1499</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>740,1319.5,740,1321.5</points>
<connection>
<GID>1022</GID>
<name>OUT</name></connection>
<intersection>1319.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>740,1319.5,740.5,1319.5</points>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection>
<intersection>740 0</intersection></hsegment></shape></wire>
<wire>
<ID>1500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>746.5,1317.5,748,1317.5</points>
<connection>
<GID>1033</GID>
<name>OUT</name></connection>
<connection>
<GID>1035</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1501</ID>
<shape>
<vsegment>
<ID>14</ID>
<points>748,1319.5,748,1322.5</points>
<connection>
<GID>1035</GID>
<name>IN_0</name></connection>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1515</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>754,1318.5,754,1318.5</points>
<connection>
<GID>1035</GID>
<name>OUT</name></connection>
<connection>
<GID>1174</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>701.5,1342,701.5,1342</points>
<connection>
<GID>1177</GID>
<name>carry_out</name></connection>
<connection>
<GID>1179</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>1519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532,1318.5,532,1318.5</points>
<connection>
<GID>1192</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1412</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1532</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>698.5,1348,698.5,1349.5</points>
<connection>
<GID>1177</GID>
<name>IN_0</name></connection>
<intersection>1349.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>698,1349.5,698.5,1349.5</points>
<connection>
<GID>1300</GID>
<name>IN_0</name></connection>
<intersection>698.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1534</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>698.5,1347,698.5,1347.5</points>
<connection>
<GID>1177</GID>
<name>IN_1</name></connection>
<intersection>1347.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>698,1347.5,698.5,1347.5</points>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection>
<intersection>698.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>1536</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>698,1345.5,698.5,1345.5</points>
<connection>
<GID>1292</GID>
<name>IN_0</name></connection>
<intersection>698.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>698.5,1345.5,698.5,1346</points>
<connection>
<GID>1177</GID>
<name>IN_2</name></connection>
<intersection>1345.5 0</intersection></vsegment></shape></wire></page 8>
<page 9>
<PageViewport>-124.789,3187.17,2293.21,1910.17</PageViewport></page 9></circuit>