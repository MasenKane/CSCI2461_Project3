<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>121.993,69.3311,197.088,31.5682</PageViewport>
<gate>
<ID>2</ID>
<type>AE_RAM_8x8</type>
<position>60.5,-4.5</position>
<input>
<ID>ADDRESS_0</ID>85 </input>
<input>
<ID>ADDRESS_1</ID>89 </input>
<input>
<ID>ADDRESS_2</ID>84 </input>
<input>
<ID>ADDRESS_3</ID>87 </input>
<input>
<ID>ADDRESS_4</ID>86 </input>
<input>
<ID>ADDRESS_5</ID>88 </input>
<input>
<ID>ADDRESS_6</ID>90 </input>
<input>
<ID>ADDRESS_7</ID>83 </input>
<input>
<ID>DATA_IN_0</ID>27 </input>
<input>
<ID>DATA_IN_1</ID>28 </input>
<input>
<ID>DATA_IN_2</ID>29 </input>
<input>
<ID>DATA_IN_3</ID>30 </input>
<input>
<ID>DATA_IN_4</ID>31 </input>
<input>
<ID>DATA_IN_5</ID>32 </input>
<input>
<ID>DATA_IN_6</ID>33 </input>
<input>
<ID>DATA_IN_7</ID>34 </input>
<output>
<ID>DATA_OUT_0</ID>27 </output>
<output>
<ID>DATA_OUT_1</ID>28 </output>
<output>
<ID>DATA_OUT_2</ID>29 </output>
<output>
<ID>DATA_OUT_3</ID>30 </output>
<output>
<ID>DATA_OUT_4</ID>31 </output>
<output>
<ID>DATA_OUT_5</ID>32 </output>
<output>
<ID>DATA_OUT_6</ID>33 </output>
<output>
<ID>DATA_OUT_7</ID>34 </output>
<input>
<ID>ENABLE_0</ID>25 </input>
<input>
<ID>write_clock</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 21</lparam>
<lparam>Address:1 21</lparam>
<lparam>Address:2 148</lparam>
<lparam>Address:3 110</lparam>
<lparam>Address:4 255</lparam></gate>
<gate>
<ID>8</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>67,-18</position>
<input>
<ID>ENABLE_0</ID>25 </input>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>29 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_4</ID>31 </input>
<input>
<ID>IN_5</ID>32 </input>
<input>
<ID>IN_6</ID>33 </input>
<input>
<ID>IN_7</ID>34 </input>
<output>
<ID>OUT_0</ID>43 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>45 </output>
<output>
<ID>OUT_3</ID>46 </output>
<output>
<ID>OUT_4</ID>47 </output>
<output>
<ID>OUT_5</ID>48 </output>
<output>
<ID>OUT_6</ID>49 </output>
<output>
<ID>OUT_7</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>14</ID>
<type>EE_VDD</type>
<position>68,-5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>BB_CLOCK</type>
<position>25,3.5</position>
<output>
<ID>CLK</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>71.5,-18</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>73.5,-18</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>75.5,-18</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>77.5,-18</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>79.5,-18</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>167.5,61</position>
<gparam>LABEL_TEXT Output 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>81.5,-18</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>83.5,-18</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>167.5,50</position>
<gparam>LABEL_TEXT Output 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>85.5,-18</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AE_REGISTER8</type>
<position>42,-5</position>
<output>
<ID>OUT_0</ID>85 </output>
<output>
<ID>OUT_1</ID>89 </output>
<output>
<ID>OUT_2</ID>84 </output>
<output>
<ID>OUT_3</ID>87 </output>
<output>
<ID>OUT_4</ID>86 </output>
<output>
<ID>OUT_5</ID>88 </output>
<output>
<ID>OUT_6</ID>90 </output>
<output>
<ID>OUT_7</ID>83 </output>
<input>
<ID>clock</ID>91 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_MUX_2x1</type>
<position>31,-13</position>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_REGISTER8</type>
<position>110.5,50</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>147 </input>
<input>
<ID>IN_6</ID>146 </input>
<input>
<ID>IN_7</ID>145 </input>
<output>
<ID>OUT_0</ID>115 </output>
<output>
<ID>OUT_1</ID>114 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>112 </output>
<output>
<ID>OUT_4</ID>111 </output>
<output>
<ID>OUT_5</ID>110 </output>
<output>
<ID>OUT_6</ID>109 </output>
<output>
<ID>OUT_7</ID>108 </output>
<input>
<ID>clock</ID>132 </input>
<input>
<ID>load</ID>155 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_REGISTER8</type>
<position>110.5,37</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>147 </input>
<input>
<ID>IN_6</ID>146 </input>
<input>
<ID>IN_7</ID>145 </input>
<output>
<ID>OUT_0</ID>131 </output>
<output>
<ID>OUT_1</ID>122 </output>
<output>
<ID>OUT_2</ID>121 </output>
<output>
<ID>OUT_3</ID>120 </output>
<output>
<ID>OUT_4</ID>119 </output>
<output>
<ID>OUT_5</ID>118 </output>
<output>
<ID>OUT_6</ID>117 </output>
<output>
<ID>OUT_7</ID>116 </output>
<input>
<ID>clock</ID>132 </input>
<input>
<ID>load</ID>156 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_MUX_4x1</type>
<position>136,87.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>108 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>92 </input>
<output>
<ID>OUT</ID>123 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_MUX_4x1</type>
<position>136,76.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>101 </input>
<input>
<ID>IN_3</ID>93 </input>
<output>
<ID>OUT</ID>124 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_MUX_4x1</type>
<position>136,65.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>102 </input>
<input>
<ID>IN_3</ID>94 </input>
<output>
<ID>OUT</ID>125 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_MUX_4x1</type>
<position>136,56</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_2</ID>103 </input>
<input>
<ID>IN_3</ID>95 </input>
<output>
<ID>OUT</ID>126 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_MUX_4x1</type>
<position>136,45</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>104 </input>
<input>
<ID>IN_3</ID>96 </input>
<output>
<ID>OUT</ID>127 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_MUX_4x1</type>
<position>136,34</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>128 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_MUX_4x1</type>
<position>136,23.5</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>114 </input>
<input>
<ID>IN_2</ID>106 </input>
<input>
<ID>IN_3</ID>98 </input>
<output>
<ID>OUT</ID>129 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_MUX_4x1</type>
<position>136,12.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>115 </input>
<input>
<ID>IN_2</ID>107 </input>
<input>
<ID>IN_3</ID>99 </input>
<output>
<ID>OUT</ID>130 </output>
<input>
<ID>SEL_0</ID>133 </input>
<input>
<ID>SEL_1</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>81</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>168,55</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>129 </input>
<input>
<ID>IN_2</ID>128 </input>
<input>
<ID>IN_3</ID>127 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>125 </input>
<input>
<ID>IN_6</ID>124 </input>
<input>
<ID>IN_7</ID>123 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>82</ID>
<type>DD_KEYPAD_HEX</type>
<position>77.5,72.5</position>
<output>
<ID>OUT_0</ID>133 </output>
<output>
<ID>OUT_1</ID>134 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>BB_CLOCK</type>
<position>99,28.5</position>
<output>
<ID>CLK</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>111.5,83.5</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>111.5,70.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>111.5,57</position>
<gparam>LABEL_TEXT R2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>111.5,44</position>
<gparam>LABEL_TEXT R3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>76,79.5</position>
<gparam>LABEL_TEXT Read 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>DD_KEYPAD_HEX</type>
<position>77.5,58.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<output>
<ID>OUT_1</ID>144 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_MUX_4x1</type>
<position>148.5,87.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>108 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>92 </input>
<output>
<ID>OUT</ID>135 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_MUX_4x1</type>
<position>148.5,76.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>101 </input>
<input>
<ID>IN_3</ID>93 </input>
<output>
<ID>OUT</ID>136 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_MUX_4x1</type>
<position>148.5,65.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>102 </input>
<input>
<ID>IN_3</ID>94 </input>
<output>
<ID>OUT</ID>137 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_MUX_4x1</type>
<position>148.5,56</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_2</ID>103 </input>
<input>
<ID>IN_3</ID>95 </input>
<output>
<ID>OUT</ID>138 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_MUX_4x1</type>
<position>148.5,45</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>104 </input>
<input>
<ID>IN_3</ID>96 </input>
<output>
<ID>OUT</ID>139 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_MUX_4x1</type>
<position>148.5,34</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>140 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_MUX_4x1</type>
<position>148.5,23.5</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>114 </input>
<input>
<ID>IN_2</ID>106 </input>
<input>
<ID>IN_3</ID>98 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_MUX_4x1</type>
<position>148.5,12.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>115 </input>
<input>
<ID>IN_2</ID>107 </input>
<input>
<ID>IN_3</ID>99 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>143 </input>
<input>
<ID>SEL_1</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>168,44</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>141 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>139 </input>
<input>
<ID>IN_4</ID>138 </input>
<input>
<ID>IN_5</ID>137 </input>
<input>
<ID>IN_6</ID>136 </input>
<input>
<ID>IN_7</ID>135 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>76,65.5</position>
<gparam>LABEL_TEXT Read 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>DD_KEYPAD_HEX</type>
<position>93.5,59</position>
<output>
<ID>OUT_0</ID>148 </output>
<output>
<ID>OUT_1</ID>147 </output>
<output>
<ID>OUT_2</ID>146 </output>
<output>
<ID>OUT_3</ID>145 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>101</ID>
<type>DD_KEYPAD_HEX</type>
<position>93.5,47</position>
<output>
<ID>OUT_0</ID>152 </output>
<output>
<ID>OUT_1</ID>151 </output>
<output>
<ID>OUT_2</ID>150 </output>
<output>
<ID>OUT_3</ID>149 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>93.5,66</position>
<gparam>LABEL_TEXT What to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>BA_DECODER_2x4</type>
<position>95.5,92</position>
<input>
<ID>ENABLE</ID>157 </input>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT_0</ID>153 </output>
<output>
<ID>OUT_1</ID>154 </output>
<output>
<ID>OUT_2</ID>155 </output>
<output>
<ID>OUT_3</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>89.5,93.5</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>87,94</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>DD_KEYPAD_HEX</type>
<position>90.5,79.5</position>
<output>
<ID>OUT_0</ID>158 </output>
<output>
<ID>OUT_1</ID>159 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>91,86.5</position>
<gparam>LABEL_TEXT Where to Write</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AE_REGISTER8</type>
<position>110.5,76.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>147 </input>
<input>
<ID>IN_6</ID>146 </input>
<input>
<ID>IN_7</ID>145 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>98 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>96 </output>
<output>
<ID>OUT_4</ID>95 </output>
<output>
<ID>OUT_5</ID>94 </output>
<output>
<ID>OUT_6</ID>93 </output>
<output>
<ID>OUT_7</ID>92 </output>
<input>
<ID>clock</ID>132 </input>
<input>
<ID>load</ID>153 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_REGISTER8</type>
<position>110.5,63.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>150 </input>
<input>
<ID>IN_3</ID>149 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>147 </input>
<input>
<ID>IN_6</ID>146 </input>
<input>
<ID>IN_7</ID>145 </input>
<output>
<ID>OUT_0</ID>107 </output>
<output>
<ID>OUT_1</ID>106 </output>
<output>
<ID>OUT_2</ID>105 </output>
<output>
<ID>OUT_3</ID>104 </output>
<output>
<ID>OUT_4</ID>103 </output>
<output>
<ID>OUT_5</ID>102 </output>
<output>
<ID>OUT_6</ID>101 </output>
<output>
<ID>OUT_7</ID>100 </output>
<input>
<ID>clock</ID>132 </input>
<input>
<ID>load</ID>154 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>121,101</position>
<gparam>LABEL_TEXT R0 - R3</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-13,67,-5</points>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-5,67,-5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-3,65.5,3.5</points>
<connection>
<GID>2</GID>
<name>write_clock</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,3.5,65.5,3.5</points>
<connection>
<GID>16</GID>
<name>CLK</name></connection>
<intersection>29 11</intersection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>29,-12,29,3.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-21.5,64,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-21.5,65,-21.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-20.5,63,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-20.5,65,-20.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-19.5,62,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-19.5,65,-19.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-18.5,61,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-18.5,65,-18.5</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-17.5,60,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_4</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_4</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-17.5,65,-17.5</points>
<connection>
<GID>8</GID>
<name>IN_4</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-16.5,59,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_5</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_5</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-16.5,65,-16.5</points>
<connection>
<GID>8</GID>
<name>IN_5</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-15.5,58,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_6</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-15.5,65,-15.5</points>
<connection>
<GID>8</GID>
<name>IN_6</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-14.5,57,-11.5</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_7</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-14.5,65,-14.5</points>
<connection>
<GID>8</GID>
<name>IN_7</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-21.5,69.5,-20</points>
<intersection>-21.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-20,84.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>84.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-21.5,69.5,-21.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-20,84.5,-18</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20.5,69.5,-20</points>
<intersection>-20.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-20,82.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>82.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-20.5,69.5,-20.5</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-20,82.5,-18</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20,69.5,-19.5</points>
<intersection>-20 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-20,80.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>80.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-19.5,69.5,-19.5</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>80.5,-20,80.5,-18</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-20,78.5,-20</points>
<intersection>69.5 3</intersection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69.5,-20,69.5,-18.5</points>
<intersection>-20 1</intersection>
<intersection>-18.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-20,78.5,-18</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>69,-18.5,69.5,-18.5</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>69.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20,69.5,-17.5</points>
<intersection>-20 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-20,76.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>76.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-17.5,69.5,-17.5</points>
<connection>
<GID>8</GID>
<name>OUT_4</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-20,76.5,-18</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20,69.5,-16.5</points>
<intersection>-20 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-16.5,69.5,-16.5</points>
<connection>
<GID>8</GID>
<name>OUT_5</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-20,74.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>74.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,-20,74.5,-18</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20,69.5,-15.5</points>
<intersection>-20 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-20,72.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>72.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-15.5,69.5,-15.5</points>
<connection>
<GID>8</GID>
<name>OUT_6</name></connection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-20,72.5,-18</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-20,69.5,-14.5</points>
<intersection>-20 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-14.5,69.5,-14.5</points>
<connection>
<GID>8</GID>
<name>OUT_7</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-20,70.5,-20</points>
<intersection>69.5 0</intersection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-20,70.5,-18</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>-20 2</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-1,55.5,-1</points>
<connection>
<GID>2</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>68</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-6,55.5,-6</points>
<connection>
<GID>2</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>68</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-8,55.5,-8</points>
<connection>
<GID>2</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-4,55.5,-4</points>
<connection>
<GID>2</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>68</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-5,55.5,-5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>68</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-3,55.5,-3</points>
<connection>
<GID>2</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>68</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-7,55.5,-7</points>
<connection>
<GID>2</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>68</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46,-2,55.5,-2</points>
<connection>
<GID>2</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>68</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-13,41,-10</points>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-13,41,-13</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,80.5,132.5,80.5</points>
<connection>
<GID>108</GID>
<name>OUT_7</name></connection>
<intersection>132.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>132.5,80.5,132.5,90.5</points>
<intersection>80.5 1</intersection>
<intersection>90.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>132.5,90.5,145.5,90.5</points>
<connection>
<GID>90</GID>
<name>IN_3</name></connection>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>132.5 4</intersection>
<intersection>144 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>144,84.5,144,90.5</points>
<intersection>84.5 8</intersection>
<intersection>90.5 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>144,84.5,145.5,84.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>144 6</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,79.5,145.5,79.5</points>
<connection>
<GID>108</GID>
<name>OUT_6</name></connection>
<connection>
<GID>91</GID>
<name>IN_3</name></connection>
<connection>
<GID>74</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,68.5,131.5,78.5</points>
<intersection>68.5 1</intersection>
<intersection>78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,68.5,145.5,68.5</points>
<connection>
<GID>92</GID>
<name>IN_3</name></connection>
<connection>
<GID>75</GID>
<name>IN_3</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,78.5,131.5,78.5</points>
<connection>
<GID>108</GID>
<name>OUT_5</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,59,131,77.5</points>
<intersection>59 1</intersection>
<intersection>77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,59,145.5,59</points>
<connection>
<GID>93</GID>
<name>IN_3</name></connection>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,77.5,131,77.5</points>
<connection>
<GID>108</GID>
<name>OUT_4</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,48,130.5,76.5</points>
<intersection>48 1</intersection>
<intersection>76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,48,145.5,48</points>
<connection>
<GID>94</GID>
<name>IN_3</name></connection>
<connection>
<GID>77</GID>
<name>IN_3</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,76.5,130.5,76.5</points>
<connection>
<GID>108</GID>
<name>OUT_3</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,37,130,75.5</points>
<intersection>37 1</intersection>
<intersection>75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,37,145.5,37</points>
<connection>
<GID>95</GID>
<name>IN_3</name></connection>
<connection>
<GID>78</GID>
<name>IN_3</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,75.5,130,75.5</points>
<connection>
<GID>108</GID>
<name>OUT_2</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,26.5,129.5,74.5</points>
<intersection>26.5 1</intersection>
<intersection>74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,26.5,145.5,26.5</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<connection>
<GID>79</GID>
<name>IN_3</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,74.5,129.5,74.5</points>
<connection>
<GID>108</GID>
<name>OUT_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,15.5,129,73.5</points>
<intersection>15.5 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,73.5,129,73.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129,15.5,145.5,15.5</points>
<connection>
<GID>97</GID>
<name>IN_3</name></connection>
<connection>
<GID>80</GID>
<name>IN_3</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,67.5,128,88.5</points>
<intersection>67.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,88.5,145.5,88.5</points>
<connection>
<GID>90</GID>
<name>IN_2</name></connection>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,67.5,128,67.5</points>
<connection>
<GID>109</GID>
<name>OUT_7</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,66.5,127.5,77.5</points>
<intersection>66.5 2</intersection>
<intersection>77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,77.5,145.5,77.5</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,66.5,127.5,66.5</points>
<connection>
<GID>109</GID>
<name>OUT_6</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,65.5,133,65.5</points>
<connection>
<GID>109</GID>
<name>OUT_5</name></connection>
<intersection>133 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133,65.5,133,66.5</points>
<connection>
<GID>75</GID>
<name>IN_2</name></connection>
<intersection>65.5 1</intersection>
<intersection>66.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>133,66.5,145.5,66.5</points>
<connection>
<GID>92</GID>
<name>IN_2</name></connection>
<intersection>133 3</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,57,127,64.5</points>
<intersection>57 1</intersection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,57,145.5,57</points>
<connection>
<GID>93</GID>
<name>IN_2</name></connection>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,64.5,127,64.5</points>
<connection>
<GID>109</GID>
<name>OUT_4</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,46,126.5,63.5</points>
<intersection>46 1</intersection>
<intersection>63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,46,145.5,46</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<connection>
<GID>77</GID>
<name>IN_2</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,63.5,126.5,63.5</points>
<connection>
<GID>109</GID>
<name>OUT_3</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,35,126,62.5</points>
<intersection>35 1</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,35,145.5,35</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<connection>
<GID>78</GID>
<name>IN_2</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,62.5,126,62.5</points>
<connection>
<GID>109</GID>
<name>OUT_2</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,24.5,125.5,61.5</points>
<intersection>24.5 2</intersection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,61.5,125.5,61.5</points>
<connection>
<GID>109</GID>
<name>OUT_1</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,24.5,145.5,24.5</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<connection>
<GID>79</GID>
<name>IN_2</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,13.5,128.5,60.5</points>
<intersection>13.5 1</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,13.5,145.5,13.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>128.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,60.5,128.5,60.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,54,124,86.5</points>
<intersection>54 2</intersection>
<intersection>86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,86.5,145.5,86.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,54,124,54</points>
<connection>
<GID>71</GID>
<name>OUT_7</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,53,123.5,75.5</points>
<intersection>53 2</intersection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,75.5,145.5,75.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,53,123.5,53</points>
<connection>
<GID>71</GID>
<name>OUT_6</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,52,123,64.5</points>
<intersection>52 2</intersection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,64.5,145.5,64.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,52,123,52</points>
<connection>
<GID>71</GID>
<name>OUT_5</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,51,122.5,55</points>
<intersection>51 2</intersection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,55,145.5,55</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,51,122.5,51</points>
<connection>
<GID>71</GID>
<name>OUT_4</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,44,122,50</points>
<intersection>44 1</intersection>
<intersection>50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,44,145.5,44</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,50,122,50</points>
<connection>
<GID>71</GID>
<name>OUT_3</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,33,121.5,49</points>
<intersection>33 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,33,145.5,33</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,49,121.5,49</points>
<connection>
<GID>71</GID>
<name>OUT_2</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,22.5,121,48</points>
<intersection>22.5 1</intersection>
<intersection>48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,22.5,145.5,22.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,48,121,48</points>
<connection>
<GID>71</GID>
<name>OUT_1</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,11.5,120.5,47</points>
<intersection>11.5 2</intersection>
<intersection>47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,47,120.5,47</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120.5,11.5,145.5,11.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,41,119.5,84.5</points>
<intersection>41 2</intersection>
<intersection>84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,84.5,133,84.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,41,119.5,41</points>
<connection>
<GID>72</GID>
<name>OUT_7</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,40,119,73.5</points>
<intersection>40 2</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,73.5,145.5,73.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,40,119,40</points>
<connection>
<GID>72</GID>
<name>OUT_6</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,39,118.5,62.5</points>
<intersection>39 2</intersection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118.5,62.5,145.5,62.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,39,118.5,39</points>
<connection>
<GID>72</GID>
<name>OUT_5</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114.5,53,145.5,53</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>114.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>114.5,38,114.5,53</points>
<connection>
<GID>72</GID>
<name>OUT_4</name></connection>
<intersection>53 1</intersection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,37,117.5,42</points>
<intersection>37 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,42,145.5,42</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,37,117.5,37</points>
<connection>
<GID>72</GID>
<name>OUT_3</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,31,117,36</points>
<intersection>31 1</intersection>
<intersection>36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,31,145.5,31</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,36,117,36</points>
<connection>
<GID>72</GID>
<name>OUT_2</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,20.5,116.5,35</points>
<intersection>20.5 1</intersection>
<intersection>35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,20.5,145.5,20.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,35,116.5,35</points>
<connection>
<GID>72</GID>
<name>OUT_1</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,59,157.5,87.5</points>
<intersection>59 2</intersection>
<intersection>87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,87.5,157.5,87.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,59,163,59</points>
<connection>
<GID>81</GID>
<name>IN_7</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,58,157.5,76.5</points>
<intersection>58 2</intersection>
<intersection>76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,76.5,157.5,76.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,58,163,58</points>
<connection>
<GID>81</GID>
<name>IN_6</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,57,157.5,65.5</points>
<intersection>57 2</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,65.5,157.5,65.5</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,57,163,57</points>
<connection>
<GID>81</GID>
<name>IN_5</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139,56,163,56</points>
<connection>
<GID>81</GID>
<name>IN_4</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,45,157.5,55</points>
<intersection>45 1</intersection>
<intersection>55 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,45,157.5,45</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,55,163,55</points>
<connection>
<GID>81</GID>
<name>IN_3</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,34,157.5,54</points>
<intersection>34 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,34,157.5,34</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,54,163,54</points>
<connection>
<GID>81</GID>
<name>IN_2</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,23.5,157.5,53</points>
<intersection>23.5 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,23.5,157.5,23.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,53,163,53</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,12.5,157.5,52</points>
<intersection>12.5 2</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,52,163,52</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,12.5,157.5,12.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,9.5,116,34</points>
<intersection>9.5 1</intersection>
<intersection>34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,9.5,145.5,9.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,34,116,34</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,28.5,106,71.5</points>
<intersection>28.5 10</intersection>
<intersection>32 8</intersection>
<intersection>45 7</intersection>
<intersection>58.5 6</intersection>
<intersection>71.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>106,71.5,109.5,71.5</points>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>106,58.5,109.5,58.5</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>106,45,109.5,45</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>106,32,109.5,32</points>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>103,28.5,106,28.5</points>
<connection>
<GID>83</GID>
<name>CLK</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,17.5,137,95.5</points>
<connection>
<GID>80</GID>
<name>SEL_0</name></connection>
<connection>
<GID>79</GID>
<name>SEL_0</name></connection>
<connection>
<GID>78</GID>
<name>SEL_0</name></connection>
<connection>
<GID>77</GID>
<name>SEL_0</name></connection>
<connection>
<GID>76</GID>
<name>SEL_0</name></connection>
<connection>
<GID>75</GID>
<name>SEL_0</name></connection>
<connection>
<GID>74</GID>
<name>SEL_0</name></connection>
<connection>
<GID>73</GID>
<name>SEL_0</name></connection>
<intersection>95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,95.5,137,95.5</points>
<intersection>83.5 2</intersection>
<intersection>137 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83.5,69.5,83.5,95.5</points>
<intersection>69.5 3</intersection>
<intersection>95.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,69.5,83.5,69.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>83.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,17.5,136,95</points>
<connection>
<GID>80</GID>
<name>SEL_1</name></connection>
<connection>
<GID>79</GID>
<name>SEL_1</name></connection>
<connection>
<GID>78</GID>
<name>SEL_1</name></connection>
<connection>
<GID>77</GID>
<name>SEL_1</name></connection>
<connection>
<GID>76</GID>
<name>SEL_1</name></connection>
<connection>
<GID>75</GID>
<name>SEL_1</name></connection>
<connection>
<GID>74</GID>
<name>SEL_1</name></connection>
<connection>
<GID>73</GID>
<name>SEL_1</name></connection>
<intersection>95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,95,136,95</points>
<intersection>83 2</intersection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>83,71.5,83,95</points>
<intersection>71.5 3</intersection>
<intersection>95 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,71.5,83,71.5</points>
<connection>
<GID>82</GID>
<name>OUT_1</name></connection>
<intersection>83 2</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,48,152,87.5</points>
<intersection>48 2</intersection>
<intersection>87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,87.5,152,87.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,48,163,48</points>
<connection>
<GID>98</GID>
<name>IN_7</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,47,152,76.5</points>
<intersection>47 2</intersection>
<intersection>76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,76.5,152,76.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,47,163,47</points>
<connection>
<GID>98</GID>
<name>IN_6</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,46,152,65.5</points>
<intersection>46 2</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,65.5,152,65.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,46,163,46</points>
<connection>
<GID>98</GID>
<name>IN_5</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,45,152,56</points>
<intersection>45 2</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,56,152,56</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,45,163,45</points>
<connection>
<GID>98</GID>
<name>IN_4</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,44,163,44</points>
<connection>
<GID>98</GID>
<name>IN_3</name></connection>
<intersection>152 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>152,44,152,45</points>
<intersection>44 1</intersection>
<intersection>45 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>151.5,45,152,45</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>152 2</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,34,152,43</points>
<intersection>34 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,34,152,34</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,43,163,43</points>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,23.5,152,42</points>
<intersection>23.5 1</intersection>
<intersection>42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151.5,23.5,152,23.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152,42,163,42</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,12.5,152,41</points>
<intersection>12.5 2</intersection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,41,163,41</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151.5,12.5,152,12.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,17.5,149.5,94</points>
<connection>
<GID>97</GID>
<name>SEL_0</name></connection>
<connection>
<GID>96</GID>
<name>SEL_0</name></connection>
<connection>
<GID>95</GID>
<name>SEL_0</name></connection>
<connection>
<GID>94</GID>
<name>SEL_0</name></connection>
<connection>
<GID>93</GID>
<name>SEL_0</name></connection>
<connection>
<GID>92</GID>
<name>SEL_0</name></connection>
<connection>
<GID>91</GID>
<name>SEL_0</name></connection>
<connection>
<GID>90</GID>
<name>SEL_0</name></connection>
<intersection>94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,94,149.5,94</points>
<intersection>84.5 2</intersection>
<intersection>149.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>84.5,55.5,84.5,94</points>
<intersection>55.5 3</intersection>
<intersection>94 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>82.5,55.5,84.5,55.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>84.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,17.5,148.5,94.5</points>
<connection>
<GID>97</GID>
<name>SEL_1</name></connection>
<connection>
<GID>96</GID>
<name>SEL_1</name></connection>
<connection>
<GID>95</GID>
<name>SEL_1</name></connection>
<connection>
<GID>94</GID>
<name>SEL_1</name></connection>
<connection>
<GID>93</GID>
<name>SEL_1</name></connection>
<connection>
<GID>92</GID>
<name>SEL_1</name></connection>
<connection>
<GID>91</GID>
<name>SEL_1</name></connection>
<connection>
<GID>90</GID>
<name>SEL_1</name></connection>
<intersection>94.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>84,94.5,148.5,94.5</points>
<intersection>84 16</intersection>
<intersection>148.5 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>84,57.5,84,94.5</points>
<intersection>57.5 18</intersection>
<intersection>94.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>82.5,57.5,84,57.5</points>
<connection>
<GID>89</GID>
<name>OUT_1</name></connection>
<intersection>84 16</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,41,105,80.5</points>
<intersection>41 6</intersection>
<intersection>54 3</intersection>
<intersection>62 4</intersection>
<intersection>67.5 2</intersection>
<intersection>80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,80.5,106.5,80.5</points>
<connection>
<GID>108</GID>
<name>IN_7</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,67.5,106.5,67.5</points>
<connection>
<GID>109</GID>
<name>IN_7</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105,54,106.5,54</points>
<connection>
<GID>71</GID>
<name>IN_7</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>98.5,62,105,62</points>
<connection>
<GID>100</GID>
<name>OUT_3</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105,41,106.5,41</points>
<connection>
<GID>72</GID>
<name>IN_7</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,40,104.5,79.5</points>
<intersection>40 6</intersection>
<intersection>53 5</intersection>
<intersection>60 2</intersection>
<intersection>66.5 3</intersection>
<intersection>79.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,60,104.5,60</points>
<connection>
<GID>100</GID>
<name>OUT_2</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,66.5,106.5,66.5</points>
<connection>
<GID>109</GID>
<name>IN_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104.5,79.5,106.5,79.5</points>
<connection>
<GID>108</GID>
<name>IN_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>104.5,53,106.5,53</points>
<connection>
<GID>71</GID>
<name>IN_6</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104.5,40,106.5,40</points>
<connection>
<GID>72</GID>
<name>IN_6</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,39,104,78.5</points>
<intersection>39 6</intersection>
<intersection>52 3</intersection>
<intersection>58 2</intersection>
<intersection>65.5 4</intersection>
<intersection>78.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,58,104,58</points>
<connection>
<GID>100</GID>
<name>OUT_1</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,52,106.5,52</points>
<connection>
<GID>71</GID>
<name>IN_5</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104,65.5,106.5,65.5</points>
<connection>
<GID>109</GID>
<name>IN_5</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>104,78.5,106.5,78.5</points>
<connection>
<GID>108</GID>
<name>IN_5</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>104,39,106.5,39</points>
<connection>
<GID>72</GID>
<name>IN_5</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,38,103.5,77.5</points>
<intersection>38 6</intersection>
<intersection>51 3</intersection>
<intersection>56 2</intersection>
<intersection>64.5 4</intersection>
<intersection>77.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,56,103.5,56</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103.5,51,106.5,51</points>
<connection>
<GID>71</GID>
<name>IN_4</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103.5,64.5,106.5,64.5</points>
<connection>
<GID>109</GID>
<name>IN_4</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103.5,77.5,106.5,77.5</points>
<connection>
<GID>108</GID>
<name>IN_4</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103.5,38,106.5,38</points>
<connection>
<GID>72</GID>
<name>IN_4</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,37,103,76.5</points>
<intersection>37 5</intersection>
<intersection>50 2</intersection>
<intersection>63.5 3</intersection>
<intersection>76.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,50,106.5,50</points>
<connection>
<GID>101</GID>
<name>OUT_3</name></connection>
<connection>
<GID>71</GID>
<name>IN_3</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>103,63.5,106.5,63.5</points>
<connection>
<GID>109</GID>
<name>IN_3</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>103,76.5,106.5,76.5</points>
<connection>
<GID>108</GID>
<name>IN_3</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,37,106.5,37</points>
<connection>
<GID>72</GID>
<name>IN_3</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,36,102.5,75.5</points>
<intersection>36 5</intersection>
<intersection>48 2</intersection>
<intersection>49 4</intersection>
<intersection>62.5 3</intersection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102.5,75.5,106.5,75.5</points>
<connection>
<GID>108</GID>
<name>IN_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,48,102.5,48</points>
<connection>
<GID>101</GID>
<name>OUT_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102.5,62.5,106.5,62.5</points>
<connection>
<GID>109</GID>
<name>IN_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102.5,49,106.5,49</points>
<connection>
<GID>71</GID>
<name>IN_2</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102.5,36,106.5,36</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,35,102,74.5</points>
<intersection>35 5</intersection>
<intersection>46 2</intersection>
<intersection>48 4</intersection>
<intersection>61.5 3</intersection>
<intersection>74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,74.5,106.5,74.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,46,102,46</points>
<connection>
<GID>101</GID>
<name>OUT_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>102,61.5,106.5,61.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102,48,106.5,48</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102,35,106.5,35</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,34,101.5,73.5</points>
<intersection>34 5</intersection>
<intersection>44 2</intersection>
<intersection>47 4</intersection>
<intersection>60.5 3</intersection>
<intersection>73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,73.5,106.5,73.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,44,101.5,44</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,60.5,106.5,60.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>101.5,47,106.5,47</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>101.5,34,106.5,34</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,82.5,108.5,90.5</points>
<intersection>82.5 2</intersection>
<intersection>90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,90.5,108.5,90.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,82.5,109.5,82.5</points>
<connection>
<GID>108</GID>
<name>load</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,69.5,108.5,91.5</points>
<intersection>69.5 2</intersection>
<intersection>91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,91.5,108.5,91.5</points>
<connection>
<GID>103</GID>
<name>OUT_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,69.5,109.5,69.5</points>
<connection>
<GID>109</GID>
<name>load</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,56,108.5,92.5</points>
<intersection>56 2</intersection>
<intersection>92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,92.5,108.5,92.5</points>
<connection>
<GID>103</GID>
<name>OUT_2</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,56,109.5,56</points>
<connection>
<GID>71</GID>
<name>load</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,43,108.5,93.5</points>
<intersection>43 2</intersection>
<intersection>93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,93.5,108.5,93.5</points>
<connection>
<GID>103</GID>
<name>OUT_3</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,43,109.5,43</points>
<connection>
<GID>72</GID>
<name>load</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,93.5,92.5,93.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,76.5,97,87.5</points>
<intersection>76.5 2</intersection>
<intersection>87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,87.5,97,87.5</points>
<intersection>92 3</intersection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,76.5,97,76.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>97 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92,87.5,92,90.5</points>
<intersection>87.5 1</intersection>
<intersection>90.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>92,90.5,92.5,90.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>92 3</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,78.5,97.5,88</points>
<intersection>78.5 2</intersection>
<intersection>88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,88,97.5,88</points>
<intersection>92.5 3</intersection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,78.5,97.5,78.5</points>
<connection>
<GID>106</GID>
<name>OUT_1</name></connection>
<intersection>97.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,88,92.5,91.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>88 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 1>
<page 2>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 2>
<page 3>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 3>
<page 4>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 4>
<page 5>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 5>
<page 6>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 6>
<page 7>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 7>
<page 8>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 8>
<page 9>
<PageViewport>-1.53459e-006,0,139.4,-70.1</PageViewport></page 9></circuit>